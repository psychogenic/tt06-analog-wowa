** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/p3_opamp.sch
.subckt p3_opamp VDD VSS PLUS MINUS VOUT
*.PININFO VDD:B VSS:B PLUS:B MINUS:B VOUT:B
XM3 VX VBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=4 m=1
XM6 VBIAS VBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=4 nf=4 m=1
XM7 VOUT VBIAS VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=7 nf=7 m=1
XR1 VBIAS VDD VSS sky130_fd_pr__res_xhigh_po_0p35 L=2.8 mult=1 m=1
XM2 V2 MINUS VX VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2.5 nf=1 m=1
XM1 V1 PLUS VX VSS sky130_fd_pr__nfet_01v8_lvt L=0.5 W=2.5 nf=1 m=1
XM4 V2 V2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=6 nf=6 m=1
XM5 V1 V2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=2 W=6 nf=6 m=1
XM8 VOUT V1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.5 W=20 nf=20 m=1
.ends
.end
