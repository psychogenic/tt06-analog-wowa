magic
tech sky130A
magscale 1 2
timestamp 1713420955
<< error_s >>
rect 16850 33440 16950 33530
rect 16850 33000 16970 33440
rect 16860 32790 16970 33000
rect 15990 32760 17080 32790
rect 15830 32680 17080 32760
rect 15830 32650 16550 32680
rect 13320 29560 13430 29670
rect 12670 29540 13430 29560
rect 12580 29450 13430 29540
rect 12580 29440 13110 29450
rect 13320 29140 13430 29450
rect 13320 28580 13460 29140
rect 13350 28420 13460 28580
<< viali >>
rect 6010 26220 6400 26280
rect 6600 26220 6990 26280
rect 7210 26220 7600 26280
rect 7820 26220 8210 26280
rect 8410 26220 8800 26280
rect 9010 26220 9400 26280
rect 9610 26220 10000 26280
<< metal1 >>
rect 5110 41349 5750 41350
rect 5110 40790 5779 41349
rect 6000 41200 6200 41400
rect 6600 41200 6800 41400
rect 7200 41200 7400 41400
rect 7800 41200 8000 41400
rect 8400 41200 8600 41400
rect 9000 41200 9200 41400
rect 9600 41200 9800 41400
rect 10200 41200 10400 41400
rect 10940 41351 11200 41430
rect 10939 41200 11200 41351
rect 5501 36108 5779 40790
rect 4762 35832 5779 36108
rect 4762 27142 5038 35832
rect 5501 35831 5779 35832
rect 10939 28000 11182 41200
rect 11493 36150 12117 36177
rect 11493 35820 11540 36150
rect 12060 35820 12117 36150
rect 11493 35783 12117 35820
rect 11544 31684 11836 35783
rect 12382 34413 12619 41419
rect 16440 40290 16640 40490
rect 20000 40380 20200 41400
rect 22000 40370 22200 41400
rect 13184 39553 14616 39926
rect 13184 36130 13557 39553
rect 13184 35830 13220 36130
rect 13530 35830 13557 36130
rect 13184 34870 13557 35830
rect 13180 34770 13557 34870
rect 13180 34670 14420 34770
rect 13180 34540 15220 34670
rect 12382 34207 14663 34413
rect 12382 34192 14220 34207
rect 12590 34190 14220 34192
rect 13770 33800 13780 34060
rect 14120 33800 14420 34060
rect 13770 33780 14420 33800
rect 12260 33570 14500 33640
rect 12260 33400 12330 33570
rect 12540 33400 14500 33570
rect 12260 33370 14500 33400
rect 11596 31660 11784 31684
rect 11480 31600 12760 31660
rect 14284 28895 14576 32966
rect 13475 28872 14576 28895
rect 13284 28649 14576 28872
rect 13475 28626 14576 28649
rect 12010 28110 12215 28272
rect 10939 27779 11910 28000
rect 10940 27770 11910 27779
rect 12010 27750 12210 28110
rect 12290 27783 12790 28018
rect 4800 26140 5000 27142
rect 10390 26803 10700 26840
rect 12010 26803 12215 27750
rect 12290 27420 12490 27783
rect 13735 27651 14066 27715
rect 12290 27000 12600 27420
rect 13730 27320 13740 27651
rect 14071 27320 14081 27651
rect 13735 26935 14066 27320
rect 10390 26558 12220 26803
rect 10390 26480 10700 26558
rect 5910 26280 10120 26300
rect 5910 26220 6010 26280
rect 6400 26220 6600 26280
rect 6990 26220 7210 26280
rect 7600 26220 7820 26280
rect 8210 26220 8410 26280
rect 8800 26220 9010 26280
rect 9400 26220 9610 26280
rect 10000 26220 10120 26280
rect 5910 26140 10120 26220
rect 14284 26140 14576 28626
rect 4800 25940 14576 26140
rect 14284 25894 14576 25940
<< via1 >>
rect 11540 35820 12060 36150
rect 13220 35830 13530 36130
rect 13780 33800 14120 34060
rect 12330 33400 12540 33570
rect 13740 27320 14071 27651
<< metal2 >>
rect 11493 36170 12117 36177
rect 11493 36150 13550 36170
rect 11493 35820 11540 36150
rect 12060 36130 13550 36150
rect 12060 35830 13220 36130
rect 13530 35830 13550 36130
rect 12060 35820 13550 35830
rect 11493 35790 13550 35820
rect 11493 35783 12117 35790
rect 13722 34070 14089 34083
rect 13722 34060 14120 34070
rect 13722 33800 13780 34060
rect 13722 33790 14120 33800
rect 12280 33570 12570 33615
rect 12280 33400 12330 33570
rect 12540 33400 12570 33570
rect 12280 31270 12570 33400
rect 13722 28040 14089 33790
rect 13720 27651 14090 28040
rect 13720 27320 13740 27651
rect 14071 27320 14090 27651
rect 13740 27310 14071 27320
use calibrated_comparator  x1
timestamp 1713420955
transform 1 0 33410 0 1 40570
box -19210 -8770 -7638 510
use r2r  x2
timestamp 1713400095
transform 1 0 7200 0 1 23800
box -2400 2370 3470 17600
use onehot2mux  x3
timestamp 1713420955
transform 0 -1 15320 1 0 28350
box -550 1780 3445 3920
<< labels >>
flabel metal1 10200 41200 10400 41400 0 FreeSans 1280 180 0 0 b7
port 7 nsew
flabel metal1 9600 41200 9800 41400 0 FreeSans 1280 180 0 0 b6
port 6 nsew
flabel metal1 9000 41200 9200 41400 0 FreeSans 1280 180 0 0 b5
port 5 nsew
flabel metal1 8400 41200 8600 41400 0 FreeSans 1280 180 0 0 b4
port 4 nsew
flabel metal1 7800 41200 8000 41400 0 FreeSans 1280 180 0 0 b3
port 3 nsew
flabel metal1 7200 41200 7400 41400 0 FreeSans 1280 180 0 0 b2
port 2 nsew
flabel metal1 6600 41200 6800 41400 0 FreeSans 1280 180 0 0 b1
port 1 nsew
flabel metal1 6000 41200 6200 41400 0 FreeSans 1280 180 0 0 b0
port 0 nsew
flabel metal1 20000 41200 20200 41400 0 FreeSans 1280 0 0 0 EN_N
port 8 nsew
flabel metal1 22000 41200 22200 41400 0 FreeSans 1280 0 0 0 COMPOUT
port 15 nsew
flabel metal1 12400 41200 12600 41400 0 FreeSans 1280 0 0 0 CAL
port 9 nsew
flabel metal1 13800 27000 14000 27200 0 FreeSans 1280 0 0 0 INPUT
port 10 nsew
flabel metal1 12400 27000 12600 27200 0 FreeSans 1280 0 0 0 EXTTHRESH
port 11 nsew
flabel metal1 16440 40290 16640 40490 0 FreeSans 1280 0 0 0 VCC
port 13 nsew
flabel metal1 4800 27200 5000 27400 0 FreeSans 1280 0 0 0 VSS
port 14 nsew
flabel metal1 11000 41230 11200 41430 0 FreeSans 1280 180 0 0 USEEXT
port 12 nsew
<< end >>
