magic
tech sky130A
magscale 1 2
timestamp 1713200672
<< viali >>
rect 1409 14569 1443 14603
rect 1961 14569 1995 14603
rect 2973 14569 3007 14603
rect 3985 14569 4019 14603
rect 4997 14569 5031 14603
rect 6009 14569 6043 14603
rect 7021 14569 7055 14603
rect 8033 14569 8067 14603
rect 9045 14569 9079 14603
rect 1593 14365 1627 14399
rect 2145 14365 2179 14399
rect 3157 14365 3191 14399
rect 4169 14365 4203 14399
rect 5181 14365 5215 14399
rect 6193 14365 6227 14399
rect 7205 14365 7239 14399
rect 8217 14365 8251 14399
rect 9229 14365 9263 14399
rect 11069 14365 11103 14399
rect 12081 14365 12115 14399
rect 13277 14365 13311 14399
rect 11253 14229 11287 14263
rect 12265 14229 12299 14263
rect 13093 14229 13127 14263
rect 3249 14025 3283 14059
rect 4721 14025 4755 14059
rect 1777 13889 1811 13923
rect 1869 13889 1903 13923
rect 2136 13889 2170 13923
rect 3341 13889 3375 13923
rect 3597 13889 3631 13923
rect 4813 13889 4847 13923
rect 5069 13889 5103 13923
rect 6929 13889 6963 13923
rect 7196 13889 7230 13923
rect 9514 13889 9548 13923
rect 10140 13889 10174 13923
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 1593 13685 1627 13719
rect 6193 13685 6227 13719
rect 8309 13685 8343 13719
rect 8401 13685 8435 13719
rect 11253 13685 11287 13719
rect 2789 13481 2823 13515
rect 7297 13481 7331 13515
rect 7573 13481 7607 13515
rect 10517 13481 10551 13515
rect 4445 13413 4479 13447
rect 5917 13345 5951 13379
rect 8401 13345 8435 13379
rect 8953 13345 8987 13379
rect 9321 13345 9355 13379
rect 11161 13345 11195 13379
rect 11345 13345 11379 13379
rect 1409 13277 1443 13311
rect 1676 13277 1710 13311
rect 4445 13277 4479 13311
rect 4583 13277 4617 13311
rect 4905 13277 4939 13311
rect 7389 13277 7423 13311
rect 7573 13277 7607 13311
rect 7974 13277 8008 13311
rect 8493 13277 8527 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9413 13277 9447 13311
rect 10333 13277 10367 13311
rect 10517 13277 10551 13311
rect 10790 13277 10824 13311
rect 11253 13277 11287 13311
rect 11529 13277 11563 13311
rect 11621 13277 11655 13311
rect 11713 13277 11747 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 6162 13209 6196 13243
rect 4721 13141 4755 13175
rect 4813 13141 4847 13175
rect 7849 13141 7883 13175
rect 8033 13141 8067 13175
rect 10609 13141 10643 13175
rect 10793 13141 10827 13175
rect 2881 12937 2915 12971
rect 3157 12937 3191 12971
rect 3433 12937 3467 12971
rect 4727 12937 4761 12971
rect 5365 12937 5399 12971
rect 5641 12937 5675 12971
rect 7205 12937 7239 12971
rect 8125 12937 8159 12971
rect 10793 12937 10827 12971
rect 3893 12869 3927 12903
rect 4813 12869 4847 12903
rect 5733 12869 5767 12903
rect 6009 12869 6043 12903
rect 6193 12869 6227 12903
rect 12081 12869 12115 12903
rect 1501 12801 1535 12835
rect 1768 12801 1802 12835
rect 2973 12801 3007 12835
rect 3065 12801 3099 12835
rect 3433 12801 3467 12835
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 4905 12801 4939 12835
rect 5365 12801 5399 12835
rect 5825 12801 5859 12835
rect 5917 12801 5951 12835
rect 6929 12801 6963 12835
rect 8309 12801 8343 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 8677 12801 8711 12835
rect 9137 12801 9171 12835
rect 9321 12801 9355 12835
rect 9413 12801 9447 12835
rect 10149 12801 10183 12835
rect 10297 12801 10331 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 10614 12801 10648 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 11989 12801 12023 12835
rect 3295 12665 3329 12699
rect 3893 12665 3927 12699
rect 5457 12597 5491 12631
rect 6193 12597 6227 12631
rect 9413 12597 9447 12631
rect 11897 12597 11931 12631
rect 1869 12393 1903 12427
rect 2697 12393 2731 12427
rect 4997 12393 5031 12427
rect 7941 12393 7975 12427
rect 10609 12393 10643 12427
rect 11069 12393 11103 12427
rect 4445 12325 4479 12359
rect 8309 12325 8343 12359
rect 8493 12257 8527 12291
rect 9137 12257 9171 12291
rect 9229 12257 9263 12291
rect 12081 12257 12115 12291
rect 2053 12189 2087 12223
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 4629 12189 4663 12223
rect 7481 12189 7515 12223
rect 7849 12189 7883 12223
rect 8125 12189 8159 12223
rect 8217 12189 8251 12223
rect 9027 12189 9061 12223
rect 9321 12189 9355 12223
rect 10057 12189 10091 12223
rect 10333 12189 10367 12223
rect 10425 12189 10459 12223
rect 11345 12189 11379 12223
rect 11529 12189 11563 12223
rect 11621 12189 11655 12223
rect 11713 12189 11747 12223
rect 4721 12121 4755 12155
rect 6561 12121 6595 12155
rect 9505 12121 9539 12155
rect 10241 12121 10275 12155
rect 10701 12121 10735 12155
rect 10885 12121 10919 12155
rect 11989 12121 12023 12155
rect 12348 12121 12382 12155
rect 4813 12053 4847 12087
rect 6837 12053 6871 12087
rect 7665 12053 7699 12087
rect 8217 12053 8251 12087
rect 13461 12053 13495 12087
rect 2145 11849 2179 11883
rect 3157 11849 3191 11883
rect 3341 11849 3375 11883
rect 3801 11849 3835 11883
rect 5457 11849 5491 11883
rect 5733 11849 5767 11883
rect 6377 11849 6411 11883
rect 9505 11849 9539 11883
rect 10977 11849 11011 11883
rect 4721 11781 4755 11815
rect 5549 11781 5583 11815
rect 9137 11781 9171 11815
rect 9413 11781 9447 11815
rect 12173 11781 12207 11815
rect 12541 11781 12575 11815
rect 12817 11781 12851 11815
rect 1961 11713 1995 11747
rect 2237 11713 2271 11747
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 3433 11713 3467 11747
rect 3985 11713 4019 11747
rect 4537 11713 4571 11747
rect 4813 11713 4847 11747
rect 4905 11713 4939 11747
rect 5365 11713 5399 11747
rect 6653 11713 6687 11747
rect 7941 11713 7975 11747
rect 8217 11713 8251 11747
rect 9321 11713 9355 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 12909 11713 12943 11747
rect 1869 11645 1903 11679
rect 2329 11645 2363 11679
rect 2605 11645 2639 11679
rect 2697 11645 2731 11679
rect 2881 11645 2915 11679
rect 3249 11645 3283 11679
rect 6536 11645 6570 11679
rect 6745 11645 6779 11679
rect 7021 11645 7055 11679
rect 8125 11645 8159 11679
rect 9689 11645 9723 11679
rect 10977 11645 11011 11679
rect 11529 11645 11563 11679
rect 11713 11645 11747 11679
rect 11989 11645 12023 11679
rect 12265 11645 12299 11679
rect 5089 11577 5123 11611
rect 5181 11577 5215 11611
rect 1685 11509 1719 11543
rect 2421 11509 2455 11543
rect 7757 11509 7791 11543
rect 8217 11509 8251 11543
rect 10517 11509 10551 11543
rect 1961 11305 1995 11339
rect 2789 11305 2823 11339
rect 4997 11305 5031 11339
rect 5549 11305 5583 11339
rect 5917 11305 5951 11339
rect 6285 11305 6319 11339
rect 6469 11305 6503 11339
rect 1869 11237 1903 11271
rect 8217 11237 8251 11271
rect 1501 11169 1535 11203
rect 3065 11169 3099 11203
rect 6101 11169 6135 11203
rect 11161 11169 11195 11203
rect 2973 11101 3007 11135
rect 3341 11101 3375 11135
rect 3433 11101 3467 11135
rect 4813 11101 4847 11135
rect 5825 11101 5859 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 6745 11101 6779 11135
rect 6929 11101 6963 11135
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 7297 11101 7331 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 8125 11101 8159 11135
rect 8309 11101 8343 11135
rect 9229 11101 9263 11135
rect 9321 11101 9355 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 10977 11101 11011 11135
rect 4445 11033 4479 11067
rect 4721 11033 4755 11067
rect 6561 11033 6595 11067
rect 3249 10965 3283 10999
rect 4629 10965 4663 10999
rect 7941 10965 7975 10999
rect 10333 10965 10367 10999
rect 10977 10965 11011 10999
rect 1961 10761 1995 10795
rect 2881 10761 2915 10795
rect 6653 10761 6687 10795
rect 10977 10761 11011 10795
rect 3049 10693 3083 10727
rect 3249 10693 3283 10727
rect 6193 10693 6227 10727
rect 8585 10693 8619 10727
rect 9045 10693 9079 10727
rect 10609 10693 10643 10727
rect 10839 10693 10873 10727
rect 2329 10625 2363 10659
rect 2421 10625 2455 10659
rect 6377 10625 6411 10659
rect 7665 10625 7699 10659
rect 7849 10625 7883 10659
rect 7941 10625 7975 10659
rect 8493 10625 8527 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 9689 10625 9723 10659
rect 10149 10625 10183 10659
rect 10333 10625 10367 10659
rect 10425 10625 10459 10659
rect 11621 10625 11655 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 12081 10625 12115 10659
rect 12173 10625 12207 10659
rect 12429 10625 12463 10659
rect 1501 10557 1535 10591
rect 2237 10557 2271 10591
rect 2513 10557 2547 10591
rect 6653 10557 6687 10591
rect 9965 10557 9999 10591
rect 1869 10489 1903 10523
rect 2053 10489 2087 10523
rect 7481 10489 7515 10523
rect 9413 10489 9447 10523
rect 12081 10489 12115 10523
rect 3065 10421 3099 10455
rect 4905 10421 4939 10455
rect 6469 10421 6503 10455
rect 8953 10421 8987 10455
rect 10793 10421 10827 10455
rect 13553 10421 13587 10455
rect 1777 10217 1811 10251
rect 3801 10217 3835 10251
rect 4445 10217 4479 10251
rect 5457 10217 5491 10251
rect 6009 10217 6043 10251
rect 6561 10217 6595 10251
rect 7113 10217 7147 10251
rect 9505 10217 9539 10251
rect 10149 10217 10183 10251
rect 10333 10217 10367 10251
rect 11897 10217 11931 10251
rect 12817 10217 12851 10251
rect 3617 10149 3651 10183
rect 6653 10149 6687 10183
rect 1961 10081 1995 10115
rect 2421 10081 2455 10115
rect 3065 10081 3099 10115
rect 5457 10081 5491 10115
rect 5917 10081 5951 10115
rect 6469 10081 6503 10115
rect 7021 10081 7055 10115
rect 9137 10081 9171 10115
rect 13093 10081 13127 10115
rect 2053 10013 2087 10047
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 4721 10013 4755 10047
rect 5549 10013 5583 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 6837 10013 6871 10047
rect 9321 10013 9355 10047
rect 9965 10013 9999 10047
rect 10149 10013 10183 10047
rect 12449 10013 12483 10047
rect 12725 10013 12759 10047
rect 12909 10013 12943 10047
rect 13185 10013 13219 10047
rect 2329 9945 2363 9979
rect 3341 9945 3375 9979
rect 3433 9945 3467 9979
rect 4077 9945 4111 9979
rect 4997 9945 5031 9979
rect 6561 9945 6595 9979
rect 7113 9945 7147 9979
rect 10425 9945 10459 9979
rect 12633 9945 12667 9979
rect 2237 9877 2271 9911
rect 3985 9877 4019 9911
rect 4629 9877 4663 9911
rect 4813 9877 4847 9911
rect 5181 9877 5215 9911
rect 5641 9877 5675 9911
rect 6101 9877 6135 9911
rect 12265 9877 12299 9911
rect 4905 9673 4939 9707
rect 9505 9673 9539 9707
rect 4997 9605 5031 9639
rect 7941 9605 7975 9639
rect 4721 9537 4755 9571
rect 5181 9537 5215 9571
rect 5365 9537 5399 9571
rect 7021 9537 7055 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 8125 9537 8159 9571
rect 8677 9537 8711 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 11621 9537 11655 9571
rect 11713 9537 11747 9571
rect 2053 9469 2087 9503
rect 4537 9469 4571 9503
rect 6929 9469 6963 9503
rect 7481 9469 7515 9503
rect 8953 9469 8987 9503
rect 9229 9469 9263 9503
rect 11897 9469 11931 9503
rect 1685 9401 1719 9435
rect 6653 9401 6687 9435
rect 7757 9401 7791 9435
rect 1593 9333 1627 9367
rect 6837 9333 6871 9367
rect 7297 9333 7331 9367
rect 7573 9333 7607 9367
rect 1777 9129 1811 9163
rect 3985 9129 4019 9163
rect 6101 9129 6135 9163
rect 6377 9129 6411 9163
rect 6745 9129 6779 9163
rect 7205 9129 7239 9163
rect 10333 9129 10367 9163
rect 4721 9061 4755 9095
rect 5457 9061 5491 9095
rect 5733 9061 5767 9095
rect 9873 9061 9907 9095
rect 1961 8993 1995 9027
rect 2053 8993 2087 9027
rect 3065 8993 3099 9027
rect 3157 8993 3191 9027
rect 7113 8993 7147 9027
rect 7757 8993 7791 9027
rect 7941 8993 7975 9027
rect 9597 8993 9631 9027
rect 10701 8993 10735 9027
rect 10885 8993 10919 9027
rect 11161 8993 11195 9027
rect 12173 8993 12207 9027
rect 2421 8925 2455 8959
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 4353 8925 4387 8959
rect 4905 8925 4939 8959
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 5631 8925 5665 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6377 8925 6411 8959
rect 6469 8925 6503 8959
rect 6929 8925 6963 8959
rect 7665 8925 7699 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9439 8925 9473 8959
rect 10241 8925 10275 8959
rect 10793 8925 10827 8959
rect 10977 8925 11011 8959
rect 2329 8857 2363 8891
rect 3985 8857 4019 8891
rect 7205 8857 7239 8891
rect 8953 8857 8987 8891
rect 9229 8857 9263 8891
rect 10149 8857 10183 8891
rect 11437 8857 11471 8891
rect 12440 8857 12474 8891
rect 2237 8789 2271 8823
rect 2881 8789 2915 8823
rect 3249 8789 3283 8823
rect 3801 8789 3835 8823
rect 7941 8789 7975 8823
rect 9689 8789 9723 8823
rect 11345 8789 11379 8823
rect 11805 8789 11839 8823
rect 13553 8789 13587 8823
rect 2053 8585 2087 8619
rect 4353 8585 4387 8619
rect 4981 8585 5015 8619
rect 5917 8585 5951 8619
rect 6561 8585 6595 8619
rect 7849 8585 7883 8619
rect 10701 8585 10735 8619
rect 12081 8585 12115 8619
rect 2697 8517 2731 8551
rect 5181 8517 5215 8551
rect 5365 8517 5399 8551
rect 5549 8517 5583 8551
rect 9321 8517 9355 8551
rect 2329 8449 2363 8483
rect 2421 8449 2455 8483
rect 3525 8449 3559 8483
rect 3617 8449 3651 8483
rect 4537 8449 4571 8483
rect 5733 8449 5767 8483
rect 6101 8449 6135 8483
rect 6745 8449 6779 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10057 8449 10091 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 12909 8449 12943 8483
rect 2237 8381 2271 8415
rect 2513 8381 2547 8415
rect 3433 8381 3467 8415
rect 3709 8381 3743 8415
rect 4721 8381 4755 8415
rect 7027 8381 7061 8415
rect 12817 8381 12851 8415
rect 3065 8313 3099 8347
rect 3249 8313 3283 8347
rect 4813 8313 4847 8347
rect 3157 8245 3191 8279
rect 4997 8245 5031 8279
rect 6929 8245 6963 8279
rect 11069 8245 11103 8279
rect 8217 8041 8251 8075
rect 8953 8041 8987 8075
rect 9689 8041 9723 8075
rect 3065 7973 3099 8007
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 3341 7837 3375 7871
rect 8125 7837 8159 7871
rect 8309 7837 8343 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 11253 7837 11287 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 1930 7769 1964 7803
rect 9873 7769 9907 7803
rect 9965 7769 9999 7803
rect 10333 7769 10367 7803
rect 11161 7769 11195 7803
rect 11529 7769 11563 7803
rect 11713 7769 11747 7803
rect 1593 7701 1627 7735
rect 3157 7701 3191 7735
rect 10057 7701 10091 7735
rect 11345 7701 11379 7735
rect 12081 7701 12115 7735
rect 5641 7497 5675 7531
rect 6929 7497 6963 7531
rect 9597 7497 9631 7531
rect 12173 7497 12207 7531
rect 2964 7429 2998 7463
rect 5304 7429 5338 7463
rect 10333 7429 10367 7463
rect 2697 7361 2731 7395
rect 5549 7361 5583 7395
rect 5917 7361 5951 7395
rect 6101 7361 6135 7395
rect 7113 7361 7147 7395
rect 7481 7361 7515 7395
rect 7941 7361 7975 7395
rect 8309 7361 8343 7395
rect 8861 7361 8895 7395
rect 9413 7361 9447 7395
rect 9873 7361 9907 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 11529 7361 11563 7395
rect 11897 7361 11931 7395
rect 12081 7361 12115 7395
rect 13297 7361 13331 7395
rect 5825 7293 5859 7327
rect 6009 7293 6043 7327
rect 7573 7293 7607 7327
rect 8677 7293 8711 7327
rect 9781 7293 9815 7327
rect 10793 7293 10827 7327
rect 13553 7293 13587 7327
rect 10333 7225 10367 7259
rect 11161 7225 11195 7259
rect 4077 7157 4111 7191
rect 4169 7157 4203 7191
rect 7113 7157 7147 7191
rect 10977 7157 11011 7191
rect 11713 7157 11747 7191
rect 12081 7157 12115 7191
rect 7481 6953 7515 6987
rect 9413 6953 9447 6987
rect 5549 6885 5583 6919
rect 7941 6885 7975 6919
rect 4905 6817 4939 6851
rect 6101 6817 6135 6851
rect 4445 6749 4479 6783
rect 4537 6749 4571 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 5917 6749 5951 6783
rect 6368 6749 6402 6783
rect 7757 6749 7791 6783
rect 8033 6749 8067 6783
rect 8953 6749 8987 6783
rect 9321 6749 9355 6783
rect 9505 6749 9539 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 11161 6749 11195 6783
rect 5825 6681 5859 6715
rect 4261 6613 4295 6647
rect 5273 6613 5307 6647
rect 8217 6613 8251 6647
rect 9137 6613 9171 6647
rect 10609 6613 10643 6647
rect 11069 6613 11103 6647
rect 4169 6409 4203 6443
rect 7757 6409 7791 6443
rect 11805 6409 11839 6443
rect 4353 6341 4387 6375
rect 10057 6341 10091 6375
rect 2145 6273 2179 6307
rect 2412 6273 2446 6307
rect 3617 6273 3651 6307
rect 3801 6273 3835 6307
rect 3893 6273 3927 6307
rect 3985 6273 4019 6307
rect 6101 6273 6135 6307
rect 6377 6273 6411 6307
rect 6644 6273 6678 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 9229 6273 9263 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 10241 6273 10275 6307
rect 10425 6273 10459 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11069 6273 11103 6307
rect 11345 6273 11379 6307
rect 12918 6273 12952 6307
rect 13185 6273 13219 6307
rect 8309 6205 8343 6239
rect 10333 6205 10367 6239
rect 11253 6205 11287 6239
rect 9597 6137 9631 6171
rect 3525 6069 3559 6103
rect 8769 6069 8803 6103
rect 9689 6069 9723 6103
rect 10057 6069 10091 6103
rect 10609 6069 10643 6103
rect 2605 5865 2639 5899
rect 4905 5865 4939 5899
rect 7205 5865 7239 5899
rect 7389 5865 7423 5899
rect 9321 5797 9355 5831
rect 12449 5797 12483 5831
rect 6377 5729 6411 5763
rect 2789 5661 2823 5695
rect 4353 5661 4387 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 6653 5661 6687 5695
rect 7297 5661 7331 5695
rect 7665 5661 7699 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 8953 5661 8987 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 12265 5661 12299 5695
rect 12461 5661 12495 5695
rect 4537 5593 4571 5627
rect 6132 5593 6166 5627
rect 9137 5593 9171 5627
rect 9597 5593 9631 5627
rect 4997 5525 5031 5559
rect 6469 5525 6503 5559
rect 7573 5525 7607 5559
rect 7941 5525 7975 5559
rect 9505 5525 9539 5559
rect 10241 5525 10275 5559
rect 11713 5525 11747 5559
rect 10819 5321 10853 5355
rect 2228 5253 2262 5287
rect 3801 5253 3835 5287
rect 9949 5253 9983 5287
rect 10149 5253 10183 5287
rect 10609 5253 10643 5287
rect 11805 5253 11839 5287
rect 1961 5185 1995 5219
rect 3617 5185 3651 5219
rect 3893 5185 3927 5219
rect 3985 5185 4019 5219
rect 4445 5185 4479 5219
rect 5733 5185 5767 5219
rect 7021 5185 7055 5219
rect 7205 5185 7239 5219
rect 7573 5185 7607 5219
rect 10425 5185 10459 5219
rect 11529 5185 11563 5219
rect 11621 5185 11655 5219
rect 11897 5185 11931 5219
rect 11989 5185 12023 5219
rect 4629 5117 4663 5151
rect 10333 5117 10367 5151
rect 12173 5117 12207 5151
rect 4169 5049 4203 5083
rect 6929 5049 6963 5083
rect 9781 5049 9815 5083
rect 10977 5049 11011 5083
rect 11805 5049 11839 5083
rect 3341 4981 3375 5015
rect 4261 4981 4295 5015
rect 5549 4981 5583 5015
rect 7389 4981 7423 5015
rect 9965 4981 9999 5015
rect 10793 4981 10827 5015
rect 12081 4981 12115 5015
rect 2421 4777 2455 4811
rect 8309 4777 8343 4811
rect 9965 4777 9999 4811
rect 13093 4777 13127 4811
rect 9321 4709 9355 4743
rect 9505 4709 9539 4743
rect 8125 4641 8159 4675
rect 8953 4641 8987 4675
rect 9781 4641 9815 4675
rect 10977 4641 11011 4675
rect 2605 4573 2639 4607
rect 4537 4573 4571 4607
rect 4813 4573 4847 4607
rect 4905 4573 4939 4607
rect 5181 4573 5215 4607
rect 5448 4573 5482 4607
rect 8033 4573 8067 4607
rect 8401 4573 8435 4607
rect 8769 4573 8803 4607
rect 9137 4573 9171 4607
rect 9413 4573 9447 4607
rect 10057 4573 10091 4607
rect 10885 4573 10919 4607
rect 11713 4573 11747 4607
rect 11980 4573 12014 4607
rect 4721 4505 4755 4539
rect 7788 4505 7822 4539
rect 10793 4505 10827 4539
rect 5089 4437 5123 4471
rect 6561 4437 6595 4471
rect 6653 4437 6687 4471
rect 8125 4437 8159 4471
rect 8585 4437 8619 4471
rect 10425 4437 10459 4471
rect 5641 4233 5675 4267
rect 8309 4233 8343 4267
rect 2145 4097 2179 4131
rect 2412 4097 2446 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 3985 4097 4019 4131
rect 4077 4097 4111 4131
rect 4537 4097 4571 4131
rect 5457 4097 5491 4131
rect 8125 4097 8159 4131
rect 8401 4097 8435 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 10609 4097 10643 4131
rect 4721 4029 4755 4063
rect 5273 4029 5307 4063
rect 10057 4029 10091 4063
rect 4261 3961 4295 3995
rect 8125 3961 8159 3995
rect 3525 3893 3559 3927
rect 4353 3893 4387 3927
rect 10793 3893 10827 3927
rect 2513 3689 2547 3723
rect 11989 3689 12023 3723
rect 13553 3689 13587 3723
rect 8493 3621 8527 3655
rect 9137 3621 9171 3655
rect 6101 3553 6135 3587
rect 10609 3553 10643 3587
rect 2697 3485 2731 3519
rect 4053 3485 4087 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 7573 3485 7607 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 8401 3485 8435 3519
rect 8677 3485 8711 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 10876 3485 10910 3519
rect 12173 3485 12207 3519
rect 4261 3417 4295 3451
rect 5181 3417 5215 3451
rect 6368 3417 6402 3451
rect 8309 3417 8343 3451
rect 8769 3417 8803 3451
rect 9321 3417 9355 3451
rect 12440 3417 12474 3451
rect 3893 3349 3927 3383
rect 4813 3349 4847 3383
rect 7481 3349 7515 3383
rect 6009 3145 6043 3179
rect 7113 3145 7147 3179
rect 9689 3145 9723 3179
rect 6745 3077 6779 3111
rect 6837 3077 6871 3111
rect 7656 3077 7690 3111
rect 2789 3009 2823 3043
rect 3056 3009 3090 3043
rect 4353 3009 4387 3043
rect 4629 3009 4663 3043
rect 4885 3009 4919 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 7389 3009 7423 3043
rect 8861 3009 8895 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 9597 3009 9631 3043
rect 10802 3009 10836 3043
rect 11069 3009 11103 3043
rect 9137 2941 9171 2975
rect 4537 2873 4571 2907
rect 4169 2805 4203 2839
rect 8769 2805 8803 2839
rect 3157 2601 3191 2635
rect 4997 2601 5031 2635
rect 6653 2601 6687 2635
rect 9045 2601 9079 2635
rect 13369 2601 13403 2635
rect 3801 2465 3835 2499
rect 4169 2465 4203 2499
rect 5365 2465 5399 2499
rect 1593 2397 1627 2431
rect 2329 2397 2363 2431
rect 3341 2397 3375 2431
rect 3617 2397 3651 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 5917 2397 5951 2431
rect 6837 2397 6871 2431
rect 7113 2397 7147 2431
rect 8309 2397 8343 2431
rect 9045 2397 9079 2431
rect 9321 2397 9355 2431
rect 9597 2397 9631 2431
rect 10149 2397 10183 2431
rect 10701 2397 10735 2431
rect 11897 2397 11931 2431
rect 13093 2397 13127 2431
rect 13553 2397 13587 2431
rect 9229 2329 9263 2363
rect 1409 2261 1443 2295
rect 2145 2261 2179 2295
rect 3433 2261 3467 2295
rect 4537 2261 4571 2295
rect 5733 2261 5767 2295
rect 6929 2261 6963 2295
rect 8125 2261 8159 2295
rect 9413 2261 9447 2295
rect 10333 2261 10367 2295
rect 10517 2261 10551 2295
rect 11713 2261 11747 2295
rect 12909 2261 12943 2295
<< metal1 >>
rect 1104 14714 13892 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13892 14714
rect 1104 14640 13892 14662
rect 842 14560 848 14612
rect 900 14600 906 14612
rect 1397 14603 1455 14609
rect 1397 14600 1409 14603
rect 900 14572 1409 14600
rect 900 14560 906 14572
rect 1397 14569 1409 14572
rect 1443 14569 1455 14603
rect 1397 14563 1455 14569
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1820 14572 1961 14600
rect 1820 14560 1826 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 1949 14563 2007 14569
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2924 14572 2973 14600
rect 2924 14560 2930 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 2961 14563 3019 14569
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 3973 14603 4031 14609
rect 3973 14600 3985 14603
rect 3936 14572 3985 14600
rect 3936 14560 3942 14572
rect 3973 14569 3985 14572
rect 4019 14569 4031 14603
rect 3973 14563 4031 14569
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 4948 14572 4997 14600
rect 4948 14560 4954 14572
rect 4985 14569 4997 14572
rect 5031 14569 5043 14603
rect 4985 14563 5043 14569
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5960 14572 6009 14600
rect 5960 14560 5966 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6972 14572 7021 14600
rect 6972 14560 6978 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7892 14572 8033 14600
rect 7892 14560 7898 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8996 14572 9045 14600
rect 8996 14560 9002 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9033 14563 9091 14569
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 4764 14436 9260 14464
rect 4764 14424 4770 14436
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 1762 14396 1768 14408
rect 1627 14368 1768 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 3050 14396 3056 14408
rect 2179 14368 3056 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3145 14399 3203 14405
rect 3145 14365 3157 14399
rect 3191 14396 3203 14399
rect 3510 14396 3516 14408
rect 3191 14368 3516 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 4154 14356 4160 14408
rect 4212 14356 4218 14408
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3694 14328 3700 14340
rect 3292 14300 3700 14328
rect 3292 14288 3298 14300
rect 3694 14288 3700 14300
rect 3752 14328 3758 14340
rect 5184 14328 5212 14359
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5684 14368 6193 14396
rect 5684 14356 5690 14368
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 7208 14328 7236 14359
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 9232 14405 9260 14436
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 7340 14368 8217 14396
rect 7340 14356 7346 14368
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 11020 14368 11069 14396
rect 11020 14356 11026 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 12032 14368 12081 14396
rect 12032 14356 12038 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13044 14368 13277 14396
rect 13044 14356 13050 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 3752 14300 5212 14328
rect 6196 14300 7236 14328
rect 3752 14288 3758 14300
rect 6196 14272 6224 14300
rect 6178 14220 6184 14272
rect 6236 14220 6242 14272
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 12250 14220 12256 14272
rect 12308 14220 12314 14272
rect 12986 14220 12992 14272
rect 13044 14260 13050 14272
rect 13081 14263 13139 14269
rect 13081 14260 13093 14263
rect 13044 14232 13093 14260
rect 13044 14220 13050 14232
rect 13081 14229 13093 14232
rect 13127 14229 13139 14263
rect 13081 14223 13139 14229
rect 1104 14170 13892 14192
rect 1104 14118 2658 14170
rect 2710 14118 2722 14170
rect 2774 14118 2786 14170
rect 2838 14118 2850 14170
rect 2902 14118 2914 14170
rect 2966 14118 2978 14170
rect 3030 14118 8658 14170
rect 8710 14118 8722 14170
rect 8774 14118 8786 14170
rect 8838 14118 8850 14170
rect 8902 14118 8914 14170
rect 8966 14118 8978 14170
rect 9030 14118 13892 14170
rect 1104 14096 13892 14118
rect 3234 14016 3240 14068
rect 3292 14016 3298 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 1578 13948 1584 14000
rect 1636 13988 1642 14000
rect 5534 13988 5540 14000
rect 1636 13960 5540 13988
rect 1636 13948 1642 13960
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1872 13929 1900 13960
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1452 13892 1777 13920
rect 1452 13880 1458 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 2124 13923 2182 13929
rect 2124 13889 2136 13923
rect 2170 13920 2182 13923
rect 2406 13920 2412 13932
rect 2170 13892 2412 13920
rect 2170 13889 2182 13892
rect 2124 13883 2182 13889
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 3344 13929 3372 13960
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 4816 13929 4844 13960
rect 5534 13948 5540 13960
rect 5592 13988 5598 14000
rect 5592 13960 6960 13988
rect 5592 13948 5598 13960
rect 3585 13923 3643 13929
rect 3585 13920 3597 13923
rect 3476 13892 3597 13920
rect 3476 13880 3482 13892
rect 3585 13889 3597 13892
rect 3631 13889 3643 13923
rect 3585 13883 3643 13889
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13889 4859 13923
rect 4801 13883 4859 13889
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 6932 13929 6960 13960
rect 5057 13923 5115 13929
rect 5057 13920 5069 13923
rect 4948 13892 5069 13920
rect 4948 13880 4954 13892
rect 5057 13889 5069 13892
rect 5103 13889 5115 13923
rect 5057 13883 5115 13889
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 7184 13923 7242 13929
rect 7184 13889 7196 13923
rect 7230 13920 7242 13923
rect 7466 13920 7472 13932
rect 7230 13892 7472 13920
rect 7230 13889 7242 13892
rect 7184 13883 7242 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 9490 13880 9496 13932
rect 9548 13929 9554 13932
rect 9548 13883 9560 13929
rect 10128 13923 10186 13929
rect 10128 13889 10140 13923
rect 10174 13920 10186 13923
rect 10410 13920 10416 13932
rect 10174 13892 10416 13920
rect 10174 13889 10186 13892
rect 10128 13883 10186 13889
rect 9548 13880 9554 13883
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 9858 13852 9864 13864
rect 9815 13824 9864 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 11790 13784 11796 13796
rect 4632 13756 4844 13784
rect 4632 13728 4660 13756
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 1670 13716 1676 13728
rect 1627 13688 1676 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 4614 13676 4620 13728
rect 4672 13676 4678 13728
rect 4816 13716 4844 13756
rect 10796 13756 11796 13784
rect 6178 13716 6184 13728
rect 4816 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8297 13719 8355 13725
rect 8297 13716 8309 13719
rect 7892 13688 8309 13716
rect 7892 13676 7898 13688
rect 8297 13685 8309 13688
rect 8343 13685 8355 13719
rect 8297 13679 8355 13685
rect 8386 13676 8392 13728
rect 8444 13676 8450 13728
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 10796 13716 10824 13756
rect 11790 13744 11796 13756
rect 11848 13744 11854 13796
rect 9456 13688 10824 13716
rect 9456 13676 9462 13688
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11241 13719 11299 13725
rect 11241 13716 11253 13719
rect 11204 13688 11253 13716
rect 11204 13676 11210 13688
rect 11241 13685 11253 13688
rect 11287 13685 11299 13719
rect 11241 13679 11299 13685
rect 1104 13626 13892 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13892 13626
rect 1104 13552 13892 13574
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 3970 13512 3976 13524
rect 2823 13484 3976 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 3970 13472 3976 13484
rect 4028 13512 4034 13524
rect 5626 13512 5632 13524
rect 4028 13484 5632 13512
rect 4028 13472 4034 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 7282 13472 7288 13524
rect 7340 13472 7346 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7524 13484 7573 13512
rect 7524 13472 7530 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7561 13475 7619 13481
rect 7668 13484 10180 13512
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 4890 13444 4896 13456
rect 4479 13416 4896 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 4448 13348 5488 13376
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1486 13308 1492 13320
rect 1443 13280 1492 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 1670 13317 1676 13320
rect 1664 13308 1676 13317
rect 1631 13280 1676 13308
rect 1664 13271 1676 13280
rect 1670 13268 1676 13271
rect 1728 13268 1734 13320
rect 3602 13268 3608 13320
rect 3660 13308 3666 13320
rect 4448 13317 4476 13348
rect 5460 13320 5488 13348
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5592 13348 5917 13376
rect 5592 13336 5598 13348
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 7668 13376 7696 13484
rect 9766 13444 9772 13456
rect 9048 13416 9772 13444
rect 5905 13339 5963 13345
rect 7392 13348 7696 13376
rect 7392 13320 7420 13348
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 8389 13379 8447 13385
rect 7892 13348 7972 13376
rect 7892 13336 7898 13348
rect 4433 13311 4491 13317
rect 4433 13308 4445 13311
rect 3660 13280 4445 13308
rect 3660 13268 3666 13280
rect 4433 13277 4445 13280
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4522 13268 4528 13320
rect 4580 13317 4586 13320
rect 4580 13311 4629 13317
rect 4580 13277 4583 13311
rect 4617 13277 4629 13311
rect 4580 13271 4629 13277
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 4982 13308 4988 13320
rect 4939 13280 4988 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 4580 13268 4586 13271
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5442 13268 5448 13320
rect 5500 13268 5506 13320
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7944 13317 7972 13348
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8435 13348 8953 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7944 13311 8020 13317
rect 7607 13280 7880 13308
rect 7944 13280 7974 13311
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 4724 13212 5120 13240
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 4724 13181 4752 13212
rect 4709 13175 4767 13181
rect 4709 13172 4721 13175
rect 3384 13144 4721 13172
rect 3384 13132 3390 13144
rect 4709 13141 4721 13144
rect 4755 13141 4767 13175
rect 4709 13135 4767 13141
rect 4798 13132 4804 13184
rect 4856 13132 4862 13184
rect 5092 13172 5120 13212
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6150 13243 6208 13249
rect 6150 13240 6162 13243
rect 5408 13212 6162 13240
rect 5408 13200 5414 13212
rect 6150 13209 6162 13212
rect 6196 13209 6208 13243
rect 6150 13203 6208 13209
rect 5902 13172 5908 13184
rect 5092 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 7852 13181 7880 13280
rect 7962 13277 7974 13280
rect 8008 13308 8020 13311
rect 8481 13311 8539 13317
rect 8008 13280 8432 13308
rect 8008 13277 8020 13280
rect 7962 13271 8020 13277
rect 8404 13240 8432 13280
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 9048 13308 9076 13416
rect 9766 13404 9772 13416
rect 9824 13404 9830 13456
rect 9309 13379 9367 13385
rect 9309 13345 9321 13379
rect 9355 13376 9367 13379
rect 9355 13348 10088 13376
rect 9355 13345 9367 13348
rect 9309 13339 9367 13345
rect 10060 13320 10088 13348
rect 8527 13280 9076 13308
rect 9125 13311 9183 13317
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 9140 13240 9168 13271
rect 8404 13212 9168 13240
rect 8496 13184 8524 13212
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 8478 13132 8484 13184
rect 8536 13132 8542 13184
rect 9232 13172 9260 13271
rect 9416 13240 9444 13271
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 10152 13308 10180 13484
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10468 13484 10517 13512
rect 10468 13472 10474 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10505 13475 10563 13481
rect 10600 13484 11744 13512
rect 10226 13404 10232 13456
rect 10284 13444 10290 13456
rect 10600 13444 10628 13484
rect 11606 13444 11612 13456
rect 10284 13416 10628 13444
rect 10704 13416 11612 13444
rect 10284 13404 10290 13416
rect 10704 13376 10732 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 10428 13348 10732 13376
rect 11149 13379 11207 13385
rect 10318 13308 10324 13320
rect 10152 13280 10324 13308
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10428 13240 10456 13348
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11195 13348 11345 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 10778 13311 10836 13317
rect 10551 13280 10640 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 9416 13212 10456 13240
rect 10226 13172 10232 13184
rect 9232 13144 10232 13172
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 10612 13181 10640 13280
rect 10778 13277 10790 13311
rect 10824 13308 10836 13311
rect 11054 13308 11060 13320
rect 10824 13280 11060 13308
rect 10824 13277 10836 13280
rect 10778 13271 10836 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 11716 13317 11744 13484
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11517 13311 11575 13317
rect 11287 13280 11376 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11348 13252 11376 13280
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11701 13311 11759 13317
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11701 13271 11759 13277
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 11330 13200 11336 13252
rect 11388 13200 11394 13252
rect 10597 13175 10655 13181
rect 10597 13141 10609 13175
rect 10643 13141 10655 13175
rect 10597 13135 10655 13141
rect 10778 13132 10784 13184
rect 10836 13132 10842 13184
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11532 13172 11560 13271
rect 11624 13184 11652 13271
rect 11808 13240 11836 13271
rect 11716 13212 11836 13240
rect 11716 13184 11744 13212
rect 11992 13184 12020 13271
rect 11204 13144 11560 13172
rect 11204 13132 11210 13144
rect 11606 13132 11612 13184
rect 11664 13132 11670 13184
rect 11698 13132 11704 13184
rect 11756 13132 11762 13184
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 1104 13082 13892 13104
rect 1104 13030 2658 13082
rect 2710 13030 2722 13082
rect 2774 13030 2786 13082
rect 2838 13030 2850 13082
rect 2902 13030 2914 13082
rect 2966 13030 2978 13082
rect 3030 13030 8658 13082
rect 8710 13030 8722 13082
rect 8774 13030 8786 13082
rect 8838 13030 8850 13082
rect 8902 13030 8914 13082
rect 8966 13030 8978 13082
rect 9030 13030 13892 13082
rect 1104 13008 13892 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 3050 12968 3056 12980
rect 2915 12940 3056 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3191 12940 3372 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3344 12912 3372 12940
rect 3418 12928 3424 12980
rect 3476 12928 3482 12980
rect 3602 12928 3608 12980
rect 3660 12928 3666 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4715 12971 4773 12977
rect 4715 12968 4727 12971
rect 4580 12940 4727 12968
rect 4580 12928 4586 12940
rect 4715 12937 4727 12940
rect 4761 12937 4773 12971
rect 4715 12931 4773 12937
rect 5350 12928 5356 12980
rect 5408 12928 5414 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 5902 12968 5908 12980
rect 5675 12940 5908 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 7374 12968 7380 12980
rect 7239 12940 7380 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 8076 12940 8125 12968
rect 8076 12928 8082 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 8113 12931 8171 12937
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10686 12968 10692 12980
rect 9824 12940 10692 12968
rect 9824 12928 9830 12940
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 10778 12928 10784 12980
rect 10836 12928 10842 12980
rect 2976 12872 3188 12900
rect 1489 12835 1547 12841
rect 1489 12801 1501 12835
rect 1535 12832 1547 12835
rect 1578 12832 1584 12844
rect 1535 12804 1584 12832
rect 1535 12801 1547 12804
rect 1489 12795 1547 12801
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 1762 12841 1768 12844
rect 1756 12795 1768 12841
rect 1762 12792 1768 12795
rect 1820 12792 1826 12844
rect 2976 12841 3004 12872
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12801 3019 12835
rect 2961 12795 3019 12801
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 3068 12628 3096 12795
rect 3160 12764 3188 12872
rect 3326 12860 3332 12912
rect 3384 12860 3390 12912
rect 3620 12900 3648 12928
rect 3528 12872 3648 12900
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12830 3479 12835
rect 3528 12830 3556 12872
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 3936 12872 4752 12900
rect 3936 12860 3942 12872
rect 4724 12844 4752 12872
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 5721 12903 5779 12909
rect 5721 12900 5733 12903
rect 4856 12872 5733 12900
rect 4856 12860 4862 12872
rect 5092 12844 5120 12872
rect 5721 12869 5733 12872
rect 5767 12900 5779 12903
rect 5997 12903 6055 12909
rect 5997 12900 6009 12903
rect 5767 12872 6009 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 5997 12869 6009 12872
rect 6043 12869 6055 12903
rect 5997 12863 6055 12869
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 7282 12900 7288 12912
rect 6236 12872 7288 12900
rect 6236 12860 6242 12872
rect 7282 12860 7288 12872
rect 7340 12860 7346 12912
rect 8404 12872 9444 12900
rect 3467 12802 3556 12830
rect 3605 12835 3663 12841
rect 3467 12801 3479 12802
rect 3421 12795 3479 12801
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3743 12804 4200 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3620 12764 3648 12795
rect 3160 12736 3648 12764
rect 3160 12708 3188 12736
rect 3142 12656 3148 12708
rect 3200 12656 3206 12708
rect 3283 12699 3341 12705
rect 3283 12665 3295 12699
rect 3329 12696 3341 12699
rect 3881 12699 3939 12705
rect 3881 12696 3893 12699
rect 3329 12668 3893 12696
rect 3329 12665 3341 12668
rect 3283 12659 3341 12665
rect 3881 12665 3893 12668
rect 3927 12665 3939 12699
rect 3881 12659 3939 12665
rect 4172 12696 4200 12804
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12832 4951 12835
rect 4939 12804 5028 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 5000 12776 5028 12804
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5353 12795 5411 12801
rect 5736 12804 5825 12832
rect 4982 12724 4988 12776
rect 5040 12724 5046 12776
rect 5368 12764 5396 12795
rect 5736 12776 5764 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 5905 12835 5963 12841
rect 5905 12832 5917 12835
rect 5859 12804 5917 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5905 12801 5917 12804
rect 5951 12801 5963 12835
rect 5905 12795 5963 12801
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 8404 12841 8432 12872
rect 9416 12844 9444 12872
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 5442 12764 5448 12776
rect 5368 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 5810 12696 5816 12708
rect 4172 12668 5816 12696
rect 4172 12628 4200 12668
rect 5810 12656 5816 12668
rect 5868 12656 5874 12708
rect 8312 12696 8340 12795
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 8662 12792 8668 12844
rect 8720 12792 8726 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 9214 12832 9220 12844
rect 9171 12804 9220 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 9324 12764 9352 12795
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 9784 12832 9812 12928
rect 11606 12900 11612 12912
rect 10336 12872 11612 12900
rect 10336 12841 10364 12872
rect 11606 12860 11612 12872
rect 11664 12900 11670 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 11664 12872 12081 12900
rect 11664 12860 11670 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 12069 12863 12127 12869
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 9784 12804 10149 12832
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10285 12835 10364 12841
rect 10285 12801 10297 12835
rect 10331 12804 10364 12835
rect 10331 12801 10343 12804
rect 10285 12795 10343 12801
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 9582 12764 9588 12776
rect 9324 12736 9588 12764
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10520 12764 10548 12795
rect 10594 12792 10600 12844
rect 10652 12841 10658 12844
rect 10652 12832 10660 12841
rect 10652 12804 10697 12832
rect 10652 12795 10660 12804
rect 10652 12792 10658 12795
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 9784 12736 10548 12764
rect 9784 12708 9812 12736
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11716 12764 11744 12795
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 11848 12804 11989 12832
rect 11848 12792 11854 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 10928 12736 11744 12764
rect 10928 12724 10934 12736
rect 9766 12696 9772 12708
rect 8312 12668 9772 12696
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 10226 12656 10232 12708
rect 10284 12696 10290 12708
rect 10410 12696 10416 12708
rect 10284 12668 10416 12696
rect 10284 12656 10290 12668
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11330 12696 11336 12708
rect 10744 12668 11336 12696
rect 10744 12656 10750 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12158 12696 12164 12708
rect 11808 12668 12164 12696
rect 3068 12600 4200 12628
rect 5445 12631 5503 12637
rect 5445 12597 5457 12631
rect 5491 12628 5503 12631
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 5491 12600 6193 12628
rect 5491 12597 5503 12600
rect 5445 12591 5503 12597
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6181 12591 6239 12597
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 10042 12628 10048 12640
rect 9447 12600 10048 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 11808 12628 11836 12668
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 10376 12600 11836 12628
rect 11885 12631 11943 12637
rect 10376 12588 10382 12600
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 11974 12628 11980 12640
rect 11931 12600 11980 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 1104 12538 13892 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13892 12538
rect 1104 12464 13892 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1820 12396 1869 12424
rect 1820 12384 1826 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 2406 12384 2412 12436
rect 2464 12424 2470 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2464 12396 2697 12424
rect 2464 12384 2470 12396
rect 2685 12393 2697 12396
rect 2731 12393 2743 12427
rect 2685 12387 2743 12393
rect 4982 12384 4988 12436
rect 5040 12384 5046 12436
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 3234 12356 3240 12368
rect 3108 12328 3240 12356
rect 3108 12316 3114 12328
rect 3234 12316 3240 12328
rect 3292 12316 3298 12368
rect 4433 12359 4491 12365
rect 4433 12325 4445 12359
rect 4479 12356 4491 12359
rect 4706 12356 4712 12368
rect 4479 12328 4712 12356
rect 4479 12325 4491 12328
rect 4433 12319 4491 12325
rect 4706 12316 4712 12328
rect 4764 12356 4770 12368
rect 5350 12356 5356 12368
rect 4764 12328 5356 12356
rect 4764 12316 4770 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 7944 12356 7972 12387
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 8720 12396 10609 12424
rect 8720 12384 8726 12396
rect 10597 12393 10609 12396
rect 10643 12424 10655 12427
rect 10778 12424 10784 12436
rect 10643 12396 10784 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11514 12424 11520 12436
rect 11112 12396 11520 12424
rect 11112 12384 11118 12396
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 8297 12359 8355 12365
rect 8297 12356 8309 12359
rect 7944 12328 8309 12356
rect 8297 12325 8309 12328
rect 8343 12356 8355 12359
rect 9306 12356 9312 12368
rect 8343 12328 9312 12356
rect 8343 12325 8355 12328
rect 8297 12319 8355 12325
rect 7484 12260 8432 12288
rect 1762 12180 1768 12232
rect 1820 12220 1826 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1820 12192 2053 12220
rect 1820 12180 1826 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2556 12192 2697 12220
rect 2556 12180 2562 12192
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3050 12220 3056 12232
rect 2915 12192 3056 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 7484 12229 7512 12260
rect 8404 12232 8432 12260
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 9122 12248 9128 12300
rect 9180 12248 9186 12300
rect 9232 12297 9260 12328
rect 9306 12316 9312 12328
rect 9364 12316 9370 12368
rect 9876 12328 12112 12356
rect 9876 12300 9904 12328
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12257 9275 12291
rect 9398 12288 9404 12300
rect 9217 12251 9275 12257
rect 9324 12260 9404 12288
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12220 4675 12223
rect 7469 12223 7527 12229
rect 4663 12192 4936 12220
rect 4663 12189 4675 12192
rect 4617 12183 4675 12189
rect 4522 12112 4528 12164
rect 4580 12152 4586 12164
rect 4709 12155 4767 12161
rect 4709 12152 4721 12155
rect 4580 12124 4721 12152
rect 4580 12112 4586 12124
rect 4709 12121 4721 12124
rect 4755 12121 4767 12155
rect 4709 12115 4767 12121
rect 4908 12096 4936 12192
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 8159 12192 8217 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8205 12189 8217 12192
rect 8251 12220 8263 12223
rect 8294 12220 8300 12232
rect 8251 12192 8300 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 6549 12155 6607 12161
rect 6549 12152 6561 12155
rect 6328 12124 6561 12152
rect 6328 12112 6334 12124
rect 6549 12121 6561 12124
rect 6595 12121 6607 12155
rect 7852 12152 7880 12183
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 8956 12223 9076 12230
rect 9324 12229 9352 12260
rect 9398 12248 9404 12260
rect 9456 12288 9462 12300
rect 9456 12260 9628 12288
rect 9456 12248 9462 12260
rect 9600 12230 9628 12260
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 12084 12297 12112 12328
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12288 12127 12291
rect 12115 12260 12204 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 9674 12230 9680 12232
rect 8956 12220 9027 12223
rect 8444 12202 9027 12220
rect 8444 12192 8984 12202
rect 8444 12180 8450 12192
rect 9015 12189 9027 12202
rect 9061 12192 9076 12223
rect 9309 12223 9367 12229
rect 9061 12189 9073 12192
rect 9015 12183 9073 12189
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9600 12202 9680 12230
rect 9646 12192 9680 12202
rect 9309 12183 9367 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10143 12192 10333 12220
rect 8478 12152 8484 12164
rect 7852 12124 8484 12152
rect 6549 12115 6607 12121
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 9499 12161 9505 12164
rect 9493 12115 9505 12161
rect 9499 12112 9505 12115
rect 9557 12112 9563 12164
rect 9766 12112 9772 12164
rect 9824 12152 9830 12164
rect 10143 12152 10171 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 11054 12220 11060 12232
rect 10459 12192 11060 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11330 12180 11336 12232
rect 11388 12180 11394 12232
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 9824 12124 10171 12152
rect 10229 12155 10287 12161
rect 9824 12112 9830 12124
rect 10229 12121 10241 12155
rect 10275 12121 10287 12155
rect 10229 12115 10287 12121
rect 4798 12044 4804 12096
rect 4856 12044 4862 12096
rect 4890 12044 4896 12096
rect 4948 12044 4954 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 5500 12056 6837 12084
rect 5500 12044 5506 12056
rect 6825 12053 6837 12056
rect 6871 12084 6883 12087
rect 7098 12084 7104 12096
rect 6871 12056 7104 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7650 12044 7656 12096
rect 7708 12044 7714 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7892 12056 8217 12084
rect 7892 12044 7898 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 10244 12084 10272 12115
rect 10594 12112 10600 12164
rect 10652 12152 10658 12164
rect 10689 12155 10747 12161
rect 10689 12152 10701 12155
rect 10652 12124 10701 12152
rect 10652 12112 10658 12124
rect 10689 12121 10701 12124
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 10410 12084 10416 12096
rect 10244 12056 10416 12084
rect 8205 12047 8263 12053
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 10888 12084 10916 12115
rect 11146 12084 11152 12096
rect 10888 12056 11152 12084
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11532 12084 11560 12183
rect 11624 12152 11652 12183
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 12176 12220 12204 12260
rect 12176 12192 12572 12220
rect 12544 12164 12572 12192
rect 11882 12152 11888 12164
rect 11624 12124 11888 12152
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 12342 12161 12348 12164
rect 11977 12155 12035 12161
rect 11977 12121 11989 12155
rect 12023 12152 12035 12155
rect 12023 12124 12296 12152
rect 12023 12121 12035 12124
rect 11977 12115 12035 12121
rect 11606 12084 11612 12096
rect 11532 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12268 12084 12296 12124
rect 12336 12115 12348 12161
rect 12342 12112 12348 12115
rect 12400 12112 12406 12164
rect 12526 12112 12532 12164
rect 12584 12112 12590 12164
rect 12434 12084 12440 12096
rect 12268 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 12952 12056 13461 12084
rect 12952 12044 12958 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 1104 11994 13892 12016
rect 1104 11942 2658 11994
rect 2710 11942 2722 11994
rect 2774 11942 2786 11994
rect 2838 11942 2850 11994
rect 2902 11942 2914 11994
rect 2966 11942 2978 11994
rect 3030 11942 8658 11994
rect 8710 11942 8722 11994
rect 8774 11942 8786 11994
rect 8838 11942 8850 11994
rect 8902 11942 8914 11994
rect 8966 11942 8978 11994
rect 9030 11942 13892 11994
rect 1104 11920 13892 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 2179 11852 2820 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 2682 11812 2688 11824
rect 1964 11784 2688 11812
rect 1964 11753 1992 11784
rect 2682 11772 2688 11784
rect 2740 11772 2746 11824
rect 2792 11756 2820 11852
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 3108 11852 3157 11880
rect 3108 11840 3114 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3510 11880 3516 11892
rect 3375 11852 3516 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3510 11840 3516 11852
rect 3568 11880 3574 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3568 11852 3801 11880
rect 3568 11840 3574 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4798 11840 4804 11892
rect 4856 11840 4862 11892
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5224 11852 5457 11880
rect 5224 11840 5230 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5718 11840 5724 11892
rect 5776 11840 5782 11892
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5868 11852 6377 11880
rect 5868 11840 5874 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 8478 11840 8484 11892
rect 8536 11840 8542 11892
rect 9490 11880 9496 11892
rect 9232 11852 9496 11880
rect 3234 11812 3240 11824
rect 2976 11784 3240 11812
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2271 11716 2728 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1636 11648 1869 11676
rect 1636 11636 1642 11648
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2700 11685 2728 11716
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 2976 11744 3004 11784
rect 3234 11772 3240 11784
rect 3292 11812 3298 11824
rect 4709 11815 4767 11821
rect 3292 11784 3832 11812
rect 3292 11772 3298 11784
rect 3804 11756 3832 11784
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4816 11812 4844 11840
rect 5537 11815 5595 11821
rect 5537 11812 5549 11815
rect 4755 11784 5549 11812
rect 4755 11781 4767 11784
rect 4709 11775 4767 11781
rect 5537 11781 5549 11784
rect 5583 11812 5595 11815
rect 5626 11812 5632 11824
rect 5583 11784 5632 11812
rect 5583 11781 5595 11784
rect 5537 11775 5595 11781
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 8496 11812 8524 11840
rect 9122 11812 9128 11824
rect 6328 11784 7420 11812
rect 6328 11772 6334 11784
rect 2884 11716 3004 11744
rect 2884 11685 2912 11716
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2372 11648 2605 11676
rect 2372 11636 2378 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11645 2927 11679
rect 2869 11639 2927 11645
rect 1670 11500 1676 11552
rect 1728 11500 1734 11552
rect 2406 11500 2412 11552
rect 2464 11500 2470 11552
rect 2608 11540 2636 11639
rect 2700 11608 2728 11639
rect 2958 11636 2964 11688
rect 3016 11676 3022 11688
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 3016 11648 3249 11676
rect 3016 11636 3022 11648
rect 3237 11645 3249 11648
rect 3283 11645 3295 11679
rect 3436 11676 3464 11707
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 4019 11716 4537 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4525 11713 4537 11716
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 3436 11648 4200 11676
rect 3237 11639 3295 11645
rect 3142 11608 3148 11620
rect 2700 11580 3148 11608
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 4172 11552 4200 11648
rect 4816 11552 4844 11707
rect 4890 11704 4896 11756
rect 4948 11704 4954 11756
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 5408 11716 6653 11744
rect 5408 11704 5414 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 4908 11676 4936 11704
rect 6546 11685 6552 11688
rect 6524 11679 6552 11685
rect 6524 11676 6536 11679
rect 4908 11648 6536 11676
rect 6524 11645 6536 11648
rect 6524 11639 6552 11645
rect 6546 11636 6552 11639
rect 6604 11636 6610 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 7006 11636 7012 11688
rect 7064 11636 7070 11688
rect 5077 11611 5135 11617
rect 5077 11577 5089 11611
rect 5123 11608 5135 11611
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 5123 11580 5181 11608
rect 5123 11577 5135 11580
rect 5077 11571 5135 11577
rect 5169 11577 5181 11580
rect 5215 11608 5227 11611
rect 6748 11608 6776 11636
rect 5215 11580 6776 11608
rect 7392 11608 7420 11784
rect 7944 11784 9128 11812
rect 7944 11753 7972 11784
rect 9122 11772 9128 11784
rect 9180 11772 9186 11824
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8386 11744 8392 11756
rect 8251 11716 8392 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8386 11704 8392 11716
rect 8444 11744 8450 11756
rect 9232 11744 9260 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10870 11880 10876 11892
rect 10192 11852 10876 11880
rect 10192 11840 10198 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11330 11880 11336 11892
rect 11011 11852 11336 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 12342 11880 12348 11892
rect 12176 11852 12348 11880
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 9674 11812 9680 11824
rect 9447 11784 9680 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 9674 11772 9680 11784
rect 9732 11812 9738 11824
rect 11146 11812 11152 11824
rect 9732 11784 11152 11812
rect 9732 11772 9738 11784
rect 11146 11772 11152 11784
rect 11204 11812 11210 11824
rect 12176 11821 12204 11852
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12161 11815 12219 11821
rect 11204 11784 11928 11812
rect 11204 11772 11210 11784
rect 8444 11716 9260 11744
rect 8444 11704 8450 11716
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 10226 11704 10232 11756
rect 10284 11744 10290 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10284 11716 10333 11744
rect 10284 11704 10290 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10502 11744 10508 11756
rect 10321 11707 10379 11713
rect 10428 11716 10508 11744
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8294 11676 8300 11688
rect 8159 11648 8300 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 9122 11608 9128 11620
rect 7392 11580 9128 11608
rect 5215 11577 5227 11580
rect 5169 11571 5227 11577
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9324 11608 9352 11704
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10428 11676 10456 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10686 11704 10692 11756
rect 10744 11704 10750 11756
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11790 11744 11796 11756
rect 11112 11716 11796 11744
rect 11112 11704 11118 11716
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11900 11753 11928 11784
rect 12161 11781 12173 11815
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 12434 11772 12440 11824
rect 12492 11772 12498 11824
rect 12529 11815 12587 11821
rect 12529 11781 12541 11815
rect 12575 11812 12587 11815
rect 12805 11815 12863 11821
rect 12805 11812 12817 11815
rect 12575 11784 12817 11812
rect 12575 11781 12587 11784
rect 12529 11775 12587 11781
rect 12805 11781 12817 11784
rect 12851 11781 12863 11815
rect 12805 11775 12863 11781
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12452 11744 12480 11772
rect 12391 11716 12480 11744
rect 12621 11747 12679 11753
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12621 11713 12633 11747
rect 12667 11713 12679 11747
rect 12894 11744 12900 11756
rect 12621 11707 12679 11713
rect 12728 11716 12900 11744
rect 9723 11648 10456 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10704 11608 10732 11704
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11011 11648 11529 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 11146 11608 11152 11620
rect 9324 11580 10645 11608
rect 10704 11580 11152 11608
rect 3510 11540 3516 11552
rect 2608 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 4154 11500 4160 11552
rect 4212 11500 4218 11552
rect 4798 11500 4804 11552
rect 4856 11500 4862 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6236 11512 7757 11540
rect 6236 11500 6242 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8205 11543 8263 11549
rect 8205 11509 8217 11543
rect 8251 11540 8263 11543
rect 9324 11540 9352 11580
rect 8251 11512 9352 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10468 11512 10517 11540
rect 10468 11500 10474 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10617 11540 10645 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 11716 11608 11744 11639
rect 11296 11580 11744 11608
rect 11992 11608 12020 11639
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 12216 11648 12265 11676
rect 12216 11636 12222 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12636 11676 12664 11707
rect 12492 11648 12664 11676
rect 12492 11636 12498 11648
rect 12728 11608 12756 11716
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 11992 11580 12756 11608
rect 11296 11568 11302 11580
rect 11698 11540 11704 11552
rect 10617 11512 11704 11540
rect 10505 11503 10563 11509
rect 11698 11500 11704 11512
rect 11756 11540 11762 11552
rect 11992 11540 12020 11580
rect 12986 11568 12992 11620
rect 13044 11568 13050 11620
rect 11756 11512 12020 11540
rect 11756 11500 11762 11512
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 13004 11540 13032 11568
rect 12216 11512 13032 11540
rect 12216 11500 12222 11512
rect 1104 11450 13892 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13892 11450
rect 1104 11376 13892 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1949 11339 2007 11345
rect 1949 11336 1961 11339
rect 1820 11308 1961 11336
rect 1820 11296 1826 11308
rect 1949 11305 1961 11308
rect 1995 11305 2007 11339
rect 1949 11299 2007 11305
rect 2406 11296 2412 11348
rect 2464 11296 2470 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2556 11308 2789 11336
rect 2556 11296 2562 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 2777 11299 2835 11305
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3234 11336 3240 11348
rect 3108 11308 3240 11336
rect 3108 11296 3114 11308
rect 3234 11296 3240 11308
rect 3292 11336 3298 11348
rect 3694 11336 3700 11348
rect 3292 11308 3700 11336
rect 3292 11296 3298 11308
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5074 11336 5080 11348
rect 5031 11308 5080 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 5626 11336 5632 11348
rect 5583 11308 5632 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 5905 11339 5963 11345
rect 5905 11305 5917 11339
rect 5951 11305 5963 11339
rect 5905 11299 5963 11305
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6362 11336 6368 11348
rect 6319 11308 6368 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11200 1547 11203
rect 1688 11200 1716 11296
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11268 1915 11271
rect 2424 11268 2452 11296
rect 1903 11240 2452 11268
rect 1903 11237 1915 11240
rect 1857 11231 1915 11237
rect 2682 11228 2688 11280
rect 2740 11268 2746 11280
rect 3326 11268 3332 11280
rect 2740 11240 3332 11268
rect 2740 11228 2746 11240
rect 3068 11209 3096 11240
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 3510 11228 3516 11280
rect 3568 11228 3574 11280
rect 5920 11268 5948 11299
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6730 11336 6736 11348
rect 6503 11308 6736 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7374 11296 7380 11348
rect 7432 11296 7438 11348
rect 7834 11296 7840 11348
rect 7892 11296 7898 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 12158 11336 12164 11348
rect 9180 11308 12164 11336
rect 9180 11296 9186 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 7392 11268 7420 11296
rect 5920 11240 7420 11268
rect 1535 11172 1716 11200
rect 3053 11203 3111 11209
rect 1535 11169 1547 11172
rect 1489 11163 1547 11169
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3528 11200 3556 11228
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 3099 11172 3133 11200
rect 3344 11172 3556 11200
rect 5736 11172 6101 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 3344 11141 3372 11172
rect 5736 11144 5764 11172
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 7852 11200 7880 11296
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 8168 11240 8217 11268
rect 8168 11228 8174 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 9490 11228 9496 11280
rect 9548 11228 9554 11280
rect 10502 11228 10508 11280
rect 10560 11268 10566 11280
rect 10560 11240 11192 11268
rect 10560 11228 10566 11240
rect 9122 11200 9128 11212
rect 6089 11163 6147 11169
rect 6748 11172 7880 11200
rect 6748 11144 6776 11172
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 1820 11104 2973 11132
rect 1820 11092 1826 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 4154 11132 4160 11144
rect 3467 11104 4160 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 2976 11064 3004 11095
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 4856 11104 5396 11132
rect 4856 11092 4862 11104
rect 3602 11064 3608 11076
rect 2976 11036 3608 11064
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4433 11067 4491 11073
rect 4433 11064 4445 11067
rect 4120 11036 4445 11064
rect 4120 11024 4126 11036
rect 4433 11033 4445 11036
rect 4479 11033 4491 11067
rect 4433 11027 4491 11033
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 4982 11064 4988 11076
rect 4755 11036 4988 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 5368 11064 5396 11104
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5951 11104 6009 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 5997 11101 6009 11104
rect 6043 11132 6055 11135
rect 6178 11132 6184 11144
rect 6043 11104 6184 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6319 11104 6684 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 6656 11076 6684 11104
rect 6730 11092 6736 11144
rect 6788 11092 6794 11144
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7190 11132 7196 11144
rect 7147 11104 7196 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 5368 11036 6561 11064
rect 6549 11033 6561 11036
rect 6595 11033 6607 11067
rect 6549 11027 6607 11033
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 7024 11064 7052 11095
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7558 11132 7564 11144
rect 7331 11104 7564 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7852 11141 7880 11172
rect 8036 11172 9128 11200
rect 8036 11141 8064 11172
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 9508 11200 9536 11228
rect 10226 11200 10232 11212
rect 9508 11172 10232 11200
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8128 11064 8156 11095
rect 6696 11036 8156 11064
rect 8312 11064 8340 11095
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8536 11104 9229 11132
rect 8536 11092 8542 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9508 11132 9536 11172
rect 10226 11160 10232 11172
rect 10284 11200 10290 11212
rect 11164 11209 11192 11240
rect 11149 11203 11207 11209
rect 10284 11172 10364 11200
rect 10284 11160 10290 11172
rect 9355 11104 9536 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10336 11141 10364 11172
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9824 11104 10149 11132
rect 9824 11092 9830 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10502 11132 10508 11144
rect 10367 11104 10508 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 9674 11064 9680 11076
rect 8312 11036 9680 11064
rect 6696 11024 6702 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10612 11064 10640 11095
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11238 11132 11244 11144
rect 11020 11104 11244 11132
rect 11020 11092 11026 11104
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11146 11064 11152 11076
rect 9784 11036 11152 11064
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3237 10999 3295 11005
rect 3237 10996 3249 10999
rect 3016 10968 3249 10996
rect 3016 10956 3022 10968
rect 3237 10965 3249 10968
rect 3283 10996 3295 10999
rect 4080 10996 4108 11024
rect 3283 10968 4108 10996
rect 3283 10965 3295 10968
rect 3237 10959 3295 10965
rect 4614 10956 4620 11008
rect 4672 10956 4678 11008
rect 7926 10956 7932 11008
rect 7984 10956 7990 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 9784 10996 9812 11036
rect 11146 11024 11152 11036
rect 11204 11064 11210 11076
rect 11514 11064 11520 11076
rect 11204 11036 11520 11064
rect 11204 11024 11210 11036
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 8168 10968 9812 10996
rect 10321 10999 10379 11005
rect 8168 10956 8174 10968
rect 10321 10965 10333 10999
rect 10367 10996 10379 10999
rect 10686 10996 10692 11008
rect 10367 10968 10692 10996
rect 10367 10965 10379 10968
rect 10321 10959 10379 10965
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 10965 10999 11023 11005
rect 10965 10965 10977 10999
rect 11011 10996 11023 10999
rect 11790 10996 11796 11008
rect 11011 10968 11796 10996
rect 11011 10965 11023 10968
rect 10965 10959 11023 10965
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 1104 10906 13892 10928
rect 1104 10854 2658 10906
rect 2710 10854 2722 10906
rect 2774 10854 2786 10906
rect 2838 10854 2850 10906
rect 2902 10854 2914 10906
rect 2966 10854 2978 10906
rect 3030 10854 8658 10906
rect 8710 10854 8722 10906
rect 8774 10854 8786 10906
rect 8838 10854 8850 10906
rect 8902 10854 8914 10906
rect 8966 10854 8978 10906
rect 9030 10854 13892 10906
rect 1104 10832 13892 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1452 10764 1961 10792
rect 1452 10752 1458 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3142 10792 3148 10804
rect 2915 10764 3148 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7006 10792 7012 10804
rect 6687 10764 7012 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7834 10752 7840 10804
rect 7892 10752 7898 10804
rect 7926 10752 7932 10804
rect 7984 10752 7990 10804
rect 8110 10752 8116 10804
rect 8168 10752 8174 10804
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 9214 10752 9220 10804
rect 9272 10752 9278 10804
rect 10318 10792 10324 10804
rect 9324 10764 10324 10792
rect 3050 10733 3056 10736
rect 3037 10727 3056 10733
rect 3037 10693 3049 10727
rect 3037 10687 3056 10693
rect 3050 10684 3056 10687
rect 3108 10684 3114 10736
rect 3237 10727 3295 10733
rect 3237 10693 3249 10727
rect 3283 10724 3295 10727
rect 4062 10724 4068 10736
rect 3283 10696 4068 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 2314 10616 2320 10668
rect 2372 10616 2378 10668
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10656 2467 10659
rect 2774 10656 2780 10668
rect 2455 10628 2780 10656
rect 2455 10625 2467 10628
rect 2409 10619 2467 10625
rect 2774 10616 2780 10628
rect 2832 10656 2838 10668
rect 3252 10656 3280 10687
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 6181 10727 6239 10733
rect 6181 10693 6193 10727
rect 6227 10724 6239 10727
rect 7852 10724 7880 10752
rect 6227 10696 7880 10724
rect 6227 10693 6239 10696
rect 6181 10687 6239 10693
rect 2832 10628 3280 10656
rect 6365 10659 6423 10665
rect 2832 10616 2838 10628
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6730 10656 6736 10668
rect 6411 10628 6736 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 1486 10548 1492 10600
rect 1544 10548 1550 10600
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 3694 10588 3700 10600
rect 2547 10560 3700 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2041 10523 2099 10529
rect 2041 10520 2053 10523
rect 1903 10492 2053 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2041 10489 2053 10492
rect 2087 10489 2099 10523
rect 2041 10483 2099 10489
rect 2240 10452 2268 10551
rect 3694 10548 3700 10560
rect 3752 10588 3758 10600
rect 3970 10588 3976 10600
rect 3752 10560 3976 10588
rect 3752 10548 3758 10560
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7558 10588 7564 10600
rect 6687 10560 7564 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 7668 10588 7696 10619
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 7944 10665 7972 10752
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7800 10628 7849 10656
rect 7800 10616 7806 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 8128 10656 8156 10752
rect 8496 10724 8524 10752
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 8496 10696 8585 10724
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8573 10687 8631 10693
rect 8864 10696 9045 10724
rect 8864 10665 8892 10696
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9033 10687 9091 10693
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 8128 10628 8493 10656
rect 7929 10619 7987 10625
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 8386 10588 8392 10600
rect 7668 10560 8392 10588
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 7469 10523 7527 10529
rect 7469 10520 7481 10523
rect 3660 10492 7481 10520
rect 3660 10480 3666 10492
rect 4724 10464 4752 10492
rect 7469 10489 7481 10492
rect 7515 10489 7527 10523
rect 7469 10483 7527 10489
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 8496 10520 8524 10619
rect 8680 10588 8708 10619
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9232 10665 9260 10752
rect 9324 10665 9352 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 10965 10795 11023 10801
rect 10560 10764 10732 10792
rect 10560 10752 10566 10764
rect 10597 10727 10655 10733
rect 9416 10696 10272 10724
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9416 10588 9444 10696
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10656 9735 10659
rect 9723 10628 10088 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 8680 10560 9444 10588
rect 9508 10588 9536 10619
rect 10060 10600 10088 10628
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9508 10560 9965 10588
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 7800 10492 8524 10520
rect 7800 10480 7806 10492
rect 9398 10480 9404 10532
rect 9456 10480 9462 10532
rect 9582 10480 9588 10532
rect 9640 10480 9646 10532
rect 10244 10520 10272 10696
rect 10597 10693 10609 10727
rect 10643 10724 10655 10727
rect 10704 10724 10732 10764
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11054 10792 11060 10804
rect 11011 10764 11060 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11974 10752 11980 10804
rect 12032 10752 12038 10804
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 10643 10696 10732 10724
rect 10827 10727 10885 10733
rect 10643 10693 10655 10696
rect 10597 10687 10655 10693
rect 10827 10693 10839 10727
rect 10873 10724 10885 10727
rect 11238 10724 11244 10736
rect 10873 10696 11244 10724
rect 10873 10693 10885 10696
rect 10827 10687 10885 10693
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11992 10724 12020 10752
rect 12544 10724 12572 10752
rect 11992 10696 12112 10724
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 10459 10628 10732 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10336 10588 10364 10619
rect 10704 10600 10732 10628
rect 11532 10628 11621 10656
rect 11532 10600 11560 10628
rect 11609 10625 11621 10628
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 12084 10665 12112 10696
rect 12176 10696 12572 10724
rect 12176 10668 12204 10696
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 10594 10588 10600 10600
rect 10336 10560 10600 10588
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10686 10548 10692 10600
rect 10744 10548 10750 10600
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 11808 10520 11836 10616
rect 10244 10492 11836 10520
rect 2314 10452 2320 10464
rect 2240 10424 2320 10452
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 4614 10452 4620 10464
rect 3099 10424 4620 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 4893 10455 4951 10461
rect 4893 10421 4905 10455
rect 4939 10452 4951 10455
rect 5534 10452 5540 10464
rect 4939 10424 5540 10452
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6457 10455 6515 10461
rect 6457 10421 6469 10455
rect 6503 10452 6515 10455
rect 6914 10452 6920 10464
rect 6503 10424 6920 10452
rect 6503 10421 6515 10424
rect 6457 10415 6515 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9600 10452 9628 10480
rect 8987 10424 9628 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10192 10424 10793 10452
rect 10192 10412 10198 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 11992 10452 12020 10619
rect 12158 10616 12164 10668
rect 12216 10616 12222 10668
rect 12417 10659 12475 10665
rect 12417 10656 12429 10659
rect 12268 10628 12429 10656
rect 12268 10588 12296 10628
rect 12417 10625 12429 10628
rect 12463 10625 12475 10659
rect 12417 10619 12475 10625
rect 12084 10560 12296 10588
rect 12084 10529 12112 10560
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 12802 10452 12808 10464
rect 11992 10424 12808 10452
rect 10781 10415 10839 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 1104 10362 13892 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13892 10362
rect 1104 10288 13892 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1765 10251 1823 10257
rect 1765 10248 1777 10251
rect 1544 10220 1777 10248
rect 1544 10208 1550 10220
rect 1765 10217 1777 10220
rect 1811 10217 1823 10251
rect 1765 10211 1823 10217
rect 2314 10208 2320 10260
rect 2372 10208 2378 10260
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3108 10220 3801 10248
rect 3108 10208 3114 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 4212 10220 4445 10248
rect 4212 10208 4218 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 5718 10248 5724 10260
rect 5491 10220 5724 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5868 10220 6009 10248
rect 5868 10208 5874 10220
rect 5997 10217 6009 10220
rect 6043 10248 6055 10251
rect 6178 10248 6184 10260
rect 6043 10220 6184 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6178 10208 6184 10220
rect 6236 10248 6242 10260
rect 6362 10248 6368 10260
rect 6236 10220 6368 10248
rect 6236 10208 6242 10220
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6512 10220 6561 10248
rect 6512 10208 6518 10220
rect 6549 10217 6561 10220
rect 6595 10248 6607 10251
rect 7101 10251 7159 10257
rect 6595 10220 7052 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 1762 10112 1768 10124
rect 1544 10084 1768 10112
rect 1544 10072 1550 10084
rect 1762 10072 1768 10084
rect 1820 10112 1826 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1820 10084 1961 10112
rect 1820 10072 1826 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 2332 10112 2360 10208
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10180 3663 10183
rect 4246 10180 4252 10192
rect 3651 10152 4252 10180
rect 3651 10149 3663 10152
rect 3605 10143 3663 10149
rect 4246 10140 4252 10152
rect 4304 10180 4310 10192
rect 4614 10180 4620 10192
rect 4304 10152 4620 10180
rect 4304 10140 4310 10152
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 5316 10152 6653 10180
rect 5316 10140 5322 10152
rect 6641 10149 6653 10152
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 2332 10084 2421 10112
rect 1949 10075 2007 10081
rect 2409 10081 2421 10084
rect 2455 10112 2467 10115
rect 3053 10115 3111 10121
rect 3053 10112 3065 10115
rect 2455 10084 3065 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 3053 10081 3065 10084
rect 3099 10081 3111 10115
rect 5276 10112 5304 10140
rect 3053 10075 3111 10081
rect 3160 10084 5304 10112
rect 5445 10115 5503 10121
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 2498 10044 2504 10056
rect 2087 10016 2504 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2317 9979 2375 9985
rect 2317 9945 2329 9979
rect 2363 9976 2375 9979
rect 2406 9976 2412 9988
rect 2363 9948 2412 9976
rect 2363 9945 2375 9948
rect 2317 9939 2375 9945
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 3160 9976 3188 10084
rect 4172 10053 4200 10084
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5491 10084 5917 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5905 10081 5917 10084
rect 5951 10112 5963 10115
rect 5951 10084 6132 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6104 10056 6132 10084
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 7024 10121 7052 10220
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7282 10248 7288 10260
rect 7147 10220 7288 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7282 10208 7288 10220
rect 7340 10248 7346 10260
rect 7650 10248 7656 10260
rect 7340 10220 7656 10248
rect 7340 10208 7346 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9456 10220 9505 10248
rect 9456 10208 9462 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 10134 10208 10140 10260
rect 10192 10208 10198 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 10594 10248 10600 10260
rect 10367 10220 10600 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11606 10208 11612 10260
rect 11664 10208 11670 10260
rect 11698 10208 11704 10260
rect 11756 10208 11762 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12158 10248 12164 10260
rect 11931 10220 12164 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 12802 10208 12808 10260
rect 12860 10208 12866 10260
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 8996 10152 9628 10180
rect 8996 10140 9002 10152
rect 6457 10115 6515 10121
rect 6457 10112 6469 10115
rect 6420 10084 6469 10112
rect 6420 10072 6426 10084
rect 6457 10081 6469 10084
rect 6503 10081 6515 10115
rect 6457 10075 6515 10081
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7466 10112 7472 10124
rect 7055 10084 7472 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8536 10084 9137 10112
rect 8536 10072 8542 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9600 10056 9628 10152
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 11624 10180 11652 10208
rect 10100 10152 11652 10180
rect 10100 10140 10106 10152
rect 11716 10112 11744 10208
rect 13538 10140 13544 10192
rect 13596 10140 13602 10192
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 9968 10084 11284 10112
rect 11716 10084 13093 10112
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4157 10047 4215 10053
rect 3283 10016 4108 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 3160 9948 3341 9976
rect 3329 9945 3341 9948
rect 3375 9945 3387 9979
rect 3329 9939 3387 9945
rect 3421 9979 3479 9985
rect 3421 9945 3433 9979
rect 3467 9976 3479 9979
rect 3602 9976 3608 9988
rect 3467 9948 3608 9976
rect 3467 9945 3479 9948
rect 3421 9939 3479 9945
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 4080 9985 4108 10016
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 4387 10016 4721 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4709 10013 4721 10016
rect 4755 10044 4767 10047
rect 5537 10047 5595 10053
rect 4755 10016 5396 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9976 4123 9979
rect 4985 9979 5043 9985
rect 4111 9948 4936 9976
rect 4111 9945 4123 9948
rect 4065 9939 4123 9945
rect 4908 9920 4936 9948
rect 4985 9945 4997 9979
rect 5031 9976 5043 9979
rect 5074 9976 5080 9988
rect 5031 9948 5080 9976
rect 5031 9945 5043 9948
rect 4985 9939 5043 9945
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5368 9920 5396 10016
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5810 10044 5816 10056
rect 5583 10016 5816 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 6012 9976 6040 10007
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10038 6331 10047
rect 6638 10044 6644 10056
rect 6380 10038 6644 10044
rect 6319 10016 6644 10038
rect 6319 10013 6408 10016
rect 6273 10010 6408 10013
rect 6273 10007 6331 10010
rect 6638 10004 6644 10016
rect 6696 10044 6702 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6696 10016 6837 10044
rect 6696 10004 6702 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 6825 10007 6883 10013
rect 7024 10016 9321 10044
rect 6549 9979 6607 9985
rect 6549 9976 6561 9979
rect 5500 9948 5764 9976
rect 6012 9948 6224 9976
rect 5500 9936 5506 9948
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 2774 9908 2780 9920
rect 2271 9880 2780 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4522 9908 4528 9920
rect 4019 9880 4528 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 4614 9868 4620 9920
rect 4672 9868 4678 9920
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 4764 9880 4813 9908
rect 4764 9868 4770 9880
rect 4801 9877 4813 9880
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 4890 9868 4896 9920
rect 4948 9908 4954 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 4948 9880 5181 9908
rect 4948 9868 4954 9880
rect 5169 9877 5181 9880
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5629 9911 5687 9917
rect 5629 9908 5641 9911
rect 5408 9880 5641 9908
rect 5408 9868 5414 9880
rect 5629 9877 5641 9880
rect 5675 9877 5687 9911
rect 5736 9908 5764 9948
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 5736 9880 6101 9908
rect 5629 9871 5687 9877
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6196 9908 6224 9948
rect 6380 9948 6561 9976
rect 6380 9908 6408 9948
rect 6549 9945 6561 9948
rect 6595 9976 6607 9979
rect 7024 9976 7052 10016
rect 9309 10013 9321 10016
rect 9355 10044 9367 10047
rect 9490 10044 9496 10056
rect 9355 10016 9496 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 9968 10053 9996 10084
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9916 10016 9965 10044
rect 9916 10004 9922 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 10226 10044 10232 10056
rect 10183 10016 10232 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 11256 9988 11284 10084
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12250 10044 12256 10056
rect 11388 10016 12256 10044
rect 11388 10004 11394 10016
rect 12250 10004 12256 10016
rect 12308 10044 12314 10056
rect 12912 10053 12940 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12308 10016 12449 10044
rect 12308 10004 12314 10016
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13556 10044 13584 10140
rect 13219 10016 13584 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 6595 9948 7052 9976
rect 7101 9979 7159 9985
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7374 9976 7380 9988
rect 7147 9948 7380 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 7374 9936 7380 9948
rect 7432 9976 7438 9988
rect 7650 9976 7656 9988
rect 7432 9948 7656 9976
rect 7432 9936 7438 9948
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 7834 9936 7840 9988
rect 7892 9976 7898 9988
rect 10410 9976 10416 9988
rect 7892 9948 10416 9976
rect 7892 9936 7898 9948
rect 10410 9936 10416 9948
rect 10468 9936 10474 9988
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11296 9948 12379 9976
rect 11296 9936 11302 9948
rect 6196 9880 6408 9908
rect 6089 9871 6147 9877
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 11422 9908 11428 9920
rect 7616 9880 11428 9908
rect 7616 9868 7622 9880
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 12253 9911 12311 9917
rect 12253 9908 12265 9911
rect 11664 9880 12265 9908
rect 11664 9868 11670 9880
rect 12253 9877 12265 9880
rect 12299 9877 12311 9911
rect 12351 9908 12379 9948
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 12621 9979 12679 9985
rect 12621 9976 12633 9979
rect 12584 9948 12633 9976
rect 12584 9936 12590 9948
rect 12621 9945 12633 9948
rect 12667 9976 12679 9979
rect 12728 9976 12756 10007
rect 12667 9948 12756 9976
rect 12667 9945 12679 9948
rect 12621 9939 12679 9945
rect 13188 9908 13216 10007
rect 12351 9880 13216 9908
rect 12253 9871 12311 9877
rect 1104 9818 13892 9840
rect 1104 9766 2658 9818
rect 2710 9766 2722 9818
rect 2774 9766 2786 9818
rect 2838 9766 2850 9818
rect 2902 9766 2914 9818
rect 2966 9766 2978 9818
rect 3030 9766 8658 9818
rect 8710 9766 8722 9818
rect 8774 9766 8786 9818
rect 8838 9766 8850 9818
rect 8902 9766 8914 9818
rect 8966 9766 8978 9818
rect 9030 9766 13892 9818
rect 1104 9744 13892 9766
rect 4522 9664 4528 9716
rect 4580 9664 4586 9716
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4672 9676 4905 9704
rect 4672 9664 4678 9676
rect 4893 9673 4905 9676
rect 4939 9704 4951 9707
rect 5166 9704 5172 9716
rect 4939 9676 5172 9704
rect 4939 9673 4951 9676
rect 4893 9667 4951 9673
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9664 5322 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6420 9676 6868 9704
rect 6420 9664 6426 9676
rect 4540 9568 4568 9664
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4540 9540 4721 9568
rect 4709 9537 4721 9540
rect 4755 9568 4767 9571
rect 5169 9571 5227 9577
rect 4755 9540 5120 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 1762 9460 1768 9512
rect 1820 9500 1826 9512
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 1820 9472 2053 9500
rect 1820 9460 1826 9472
rect 2041 9469 2053 9472
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4890 9500 4896 9512
rect 4571 9472 4896 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5092 9500 5120 9540
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5276 9568 5304 9664
rect 6840 9636 6868 9676
rect 9490 9664 9496 9716
rect 9548 9664 9554 9716
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 11146 9704 11152 9716
rect 9640 9676 11152 9704
rect 9640 9664 9646 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 12342 9704 12348 9716
rect 11572 9676 12348 9704
rect 11572 9664 11578 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 6840 9608 7420 9636
rect 5215 9540 5304 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6840 9568 6868 9608
rect 7392 9580 7420 9608
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 7929 9639 7987 9645
rect 7929 9636 7941 9639
rect 7800 9608 7941 9636
rect 7800 9596 7806 9608
rect 7929 9605 7941 9608
rect 7975 9605 7987 9639
rect 10134 9636 10140 9648
rect 7929 9599 7987 9605
rect 9232 9608 9444 9636
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6840 9540 7021 9568
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7098 9528 7104 9580
rect 7156 9528 7162 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 7248 9540 7297 9568
rect 7248 9528 7254 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 5442 9500 5448 9512
rect 5092 9472 5448 9500
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 1670 9392 1676 9444
rect 1728 9392 1734 9444
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 6454 9432 6460 9444
rect 5132 9404 6460 9432
rect 5132 9392 5138 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6604 9404 6653 9432
rect 6604 9392 6610 9404
rect 6641 9401 6653 9404
rect 6687 9401 6699 9435
rect 6641 9395 6699 9401
rect 1578 9324 1584 9376
rect 1636 9324 1642 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 5902 9364 5908 9376
rect 3200 9336 5908 9364
rect 3200 9324 3206 9336
rect 5902 9324 5908 9336
rect 5960 9364 5966 9376
rect 6270 9364 6276 9376
rect 5960 9336 6276 9364
rect 5960 9324 5966 9336
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6748 9364 6776 9528
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 6932 9432 6960 9463
rect 7190 9432 7196 9444
rect 6932 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7300 9432 7328 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7760 9540 8125 9568
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 7558 9500 7564 9512
rect 7515 9472 7564 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7760 9441 7788 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8711 9540 9137 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 9125 9537 9137 9540
rect 9171 9568 9183 9571
rect 9232 9568 9260 9608
rect 9171 9540 9260 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 7745 9435 7803 9441
rect 7745 9432 7757 9435
rect 7300 9404 7757 9432
rect 7745 9401 7757 9404
rect 7791 9401 7803 9435
rect 8956 9432 8984 9463
rect 9030 9460 9036 9512
rect 9088 9500 9094 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9088 9472 9229 9500
rect 9088 9460 9094 9472
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9416 9500 9444 9608
rect 9508 9608 10140 9636
rect 9508 9577 9536 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 10796 9608 11744 9636
rect 10796 9580 10824 9608
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9858 9568 9864 9580
rect 9723 9540 9864 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11606 9568 11612 9580
rect 11112 9540 11612 9568
rect 11112 9528 11118 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11716 9577 11744 9608
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 9416 9472 11897 9500
rect 9217 9463 9275 9469
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 9306 9432 9312 9444
rect 8956 9404 9312 9432
rect 7745 9395 7803 9401
rect 9306 9392 9312 9404
rect 9364 9432 9370 9444
rect 11900 9432 11928 9463
rect 12526 9432 12532 9444
rect 9364 9404 9904 9432
rect 11900 9404 12532 9432
rect 9364 9392 9370 9404
rect 6822 9364 6828 9376
rect 6748 9336 6828 9364
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6972 9336 7297 9364
rect 6972 9324 6978 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 7650 9364 7656 9376
rect 7607 9336 7656 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7650 9324 7656 9336
rect 7708 9364 7714 9376
rect 9766 9364 9772 9376
rect 7708 9336 9772 9364
rect 7708 9324 7714 9336
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9876 9364 9904 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 11974 9364 11980 9376
rect 9876 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 1104 9274 13892 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13892 9274
rect 1104 9200 13892 9222
rect 1762 9120 1768 9172
rect 1820 9120 1826 9172
rect 2498 9160 2504 9172
rect 2056 9132 2504 9160
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 2056 9033 2084 9132
rect 2498 9120 2504 9132
rect 2556 9160 2562 9172
rect 3142 9160 3148 9172
rect 2556 9132 3148 9160
rect 2556 9120 2562 9132
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4246 9160 4252 9172
rect 4019 9132 4252 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5408 9132 5764 9160
rect 5408 9120 5414 9132
rect 2148 9064 3096 9092
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1544 8996 1961 9024
rect 1544 8984 1550 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2041 9027 2099 9033
rect 2041 8993 2053 9027
rect 2087 8993 2099 9027
rect 2041 8987 2099 8993
rect 1964 8956 1992 8987
rect 2148 8956 2176 9064
rect 2958 9024 2964 9036
rect 2332 8996 2964 9024
rect 2332 8956 2360 8996
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3068 9033 3096 9064
rect 3160 9033 3188 9120
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4709 9095 4767 9101
rect 4709 9092 4721 9095
rect 4120 9064 4721 9092
rect 4120 9052 4126 9064
rect 4709 9061 4721 9064
rect 4755 9061 4767 9095
rect 4709 9055 4767 9061
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5445 9095 5503 9101
rect 5445 9092 5457 9095
rect 5040 9064 5457 9092
rect 5040 9052 5046 9064
rect 5445 9061 5457 9064
rect 5491 9061 5503 9095
rect 5445 9055 5503 9061
rect 5626 9052 5632 9104
rect 5684 9052 5690 9104
rect 5736 9101 5764 9132
rect 6012 9132 6101 9160
rect 5721 9095 5779 9101
rect 5721 9061 5733 9095
rect 5767 9061 5779 9095
rect 5721 9055 5779 9061
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 8993 3111 9027
rect 3053 8987 3111 8993
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 1964 8928 2176 8956
rect 2240 8928 2360 8956
rect 2240 8829 2268 8928
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 2464 8928 3433 8956
rect 2464 8916 2470 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 3510 8916 3516 8968
rect 3568 8916 3574 8968
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4890 8956 4896 8968
rect 4387 8928 4896 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5644 8965 5672 9052
rect 6012 9024 6040 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 6362 9120 6368 9172
rect 6420 9120 6426 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6696 9132 6745 9160
rect 6696 9120 6702 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 10318 9160 10324 9172
rect 7248 9132 9674 9160
rect 7248 9120 7254 9132
rect 5920 8996 6040 9024
rect 5619 8959 5677 8965
rect 5408 8928 5488 8956
rect 5408 8916 5414 8928
rect 2314 8848 2320 8900
rect 2372 8888 2378 8900
rect 3973 8891 4031 8897
rect 2372 8860 3832 8888
rect 2372 8848 2378 8860
rect 2225 8823 2283 8829
rect 2225 8789 2237 8823
rect 2271 8789 2283 8823
rect 2225 8783 2283 8789
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2556 8792 2881 8820
rect 2556 8780 2562 8792
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3804 8829 3832 8860
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 4706 8888 4712 8900
rect 4019 8860 4712 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3108 8792 3249 8820
rect 3108 8780 3114 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8789 3847 8823
rect 5460 8820 5488 8928
rect 5619 8925 5631 8959
rect 5665 8925 5677 8959
rect 5619 8919 5677 8925
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 5920 8965 5948 8996
rect 6270 8984 6276 9036
rect 6328 8984 6334 9036
rect 6380 9024 6408 9120
rect 9490 9092 9496 9104
rect 7944 9064 9496 9092
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6380 8996 7113 9024
rect 7101 8993 7113 8996
rect 7147 9024 7159 9027
rect 7282 9024 7288 9036
rect 7147 8996 7288 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7944 9033 7972 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 9646 9092 9674 9132
rect 10152 9132 10324 9160
rect 9646 9064 9812 9092
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7432 8996 7757 9024
rect 7432 8984 7438 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 9585 9027 9643 9033
rect 9585 9006 9597 9027
rect 9631 9006 9643 9027
rect 9784 9024 9812 9064
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 10152 9092 10180 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11882 9160 11888 9172
rect 11204 9132 11888 9160
rect 11204 9120 11210 9132
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 9916 9064 10180 9092
rect 9916 9052 9922 9064
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10284 9064 10732 9092
rect 10284 9052 10290 9064
rect 10704 9033 10732 9064
rect 10689 9027 10747 9033
rect 7929 8987 7987 8993
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 6295 8956 6323 8984
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6295 8928 6377 8956
rect 5905 8919 5963 8925
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 5920 8888 5948 8919
rect 5776 8860 5948 8888
rect 6472 8888 6500 8919
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6788 8928 6929 8956
rect 6788 8916 6794 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 7650 8956 7656 8968
rect 6917 8919 6975 8925
rect 7024 8928 7656 8956
rect 7024 8888 7052 8928
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9214 8926 9220 8978
rect 9272 8956 9278 8978
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 9272 8928 9321 8956
rect 9272 8926 9278 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9427 8959 9485 8965
rect 9427 8925 9439 8959
rect 9473 8956 9485 8959
rect 9473 8928 9545 8956
rect 9582 8954 9588 9006
rect 9640 8954 9646 9006
rect 9784 8996 10456 9024
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9473 8925 9485 8928
rect 9427 8919 9485 8925
rect 6472 8860 7052 8888
rect 5776 8848 5782 8860
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7558 8888 7564 8900
rect 7248 8860 7564 8888
rect 7248 8848 7254 8860
rect 7558 8848 7564 8860
rect 7616 8888 7622 8900
rect 8588 8888 8616 8916
rect 7616 8860 8616 8888
rect 7616 8848 7622 8860
rect 8938 8848 8944 8900
rect 8996 8848 9002 8900
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 9140 8860 9229 8888
rect 9140 8832 9168 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 9517 8888 9545 8928
rect 10152 8928 10241 8956
rect 10152 8900 10180 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 9582 8888 9588 8900
rect 9517 8860 9588 8888
rect 9217 8851 9275 8857
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 10134 8848 10140 8900
rect 10192 8848 10198 8900
rect 10428 8888 10456 8996
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10873 9027 10931 9033
rect 10735 8996 10824 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10796 8965 10824 8996
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10919 8996 11161 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 12124 8996 12173 9024
rect 12124 8984 12130 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 10686 8888 10692 8900
rect 10428 8860 10692 8888
rect 10686 8848 10692 8860
rect 10744 8888 10750 8900
rect 10980 8888 11008 8919
rect 12434 8897 12440 8900
rect 11425 8891 11483 8897
rect 11425 8888 11437 8891
rect 10744 8860 11008 8888
rect 11072 8860 11437 8888
rect 10744 8848 10750 8860
rect 6822 8820 6828 8832
rect 5460 8792 6828 8820
rect 3789 8783 3847 8789
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7800 8792 7941 8820
rect 7800 8780 7806 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 9122 8780 9128 8832
rect 9180 8780 9186 8832
rect 9490 8780 9496 8832
rect 9548 8820 9554 8832
rect 9677 8823 9735 8829
rect 9677 8820 9689 8823
rect 9548 8792 9689 8820
rect 9548 8780 9554 8792
rect 9677 8789 9689 8792
rect 9723 8789 9735 8823
rect 9677 8783 9735 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 10778 8820 10784 8832
rect 9916 8792 10784 8820
rect 9916 8780 9922 8792
rect 10778 8780 10784 8792
rect 10836 8820 10842 8832
rect 11072 8820 11100 8860
rect 11425 8857 11437 8860
rect 11471 8857 11483 8891
rect 11425 8851 11483 8857
rect 12428 8851 12440 8897
rect 12434 8848 12440 8851
rect 12492 8848 12498 8900
rect 10836 8792 11100 8820
rect 11333 8823 11391 8829
rect 10836 8780 10842 8792
rect 11333 8789 11345 8823
rect 11379 8820 11391 8823
rect 11698 8820 11704 8832
rect 11379 8792 11704 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 11974 8820 11980 8832
rect 11839 8792 11980 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 1104 8730 13892 8752
rect 1104 8678 2658 8730
rect 2710 8678 2722 8730
rect 2774 8678 2786 8730
rect 2838 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 8658 8730
rect 8710 8678 8722 8730
rect 8774 8678 8786 8730
rect 8838 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 13892 8730
rect 1104 8656 13892 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2041 8619 2099 8625
rect 2041 8616 2053 8619
rect 1728 8588 2053 8616
rect 1728 8576 1734 8588
rect 2041 8585 2053 8588
rect 2087 8585 2099 8619
rect 2041 8579 2099 8585
rect 2314 8576 2320 8628
rect 2372 8576 2378 8628
rect 2498 8576 2504 8628
rect 2556 8576 2562 8628
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3108 8588 3648 8616
rect 3108 8576 3114 8588
rect 2332 8489 2360 8576
rect 2516 8548 2544 8576
rect 2685 8551 2743 8557
rect 2685 8548 2697 8551
rect 2516 8520 2697 8548
rect 2685 8517 2697 8520
rect 2731 8517 2743 8551
rect 3068 8548 3096 8576
rect 2685 8511 2743 8517
rect 2792 8520 3096 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2792 8480 2820 8520
rect 3620 8489 3648 8588
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4982 8625 4988 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4304 8588 4353 8616
rect 4304 8576 4310 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 4969 8619 4988 8625
rect 4969 8585 4981 8619
rect 4969 8579 4988 8585
rect 4982 8576 4988 8579
rect 5040 8576 5046 8628
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5902 8576 5908 8628
rect 5960 8576 5966 8628
rect 6362 8576 6368 8628
rect 6420 8576 6426 8628
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 6822 8616 6828 8628
rect 6595 8588 6828 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 10226 8616 10232 8628
rect 7944 8588 10232 8616
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 3513 8483 3571 8489
rect 3513 8480 3525 8483
rect 2455 8452 2820 8480
rect 2884 8452 3525 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 2774 8412 2780 8424
rect 2547 8384 2780 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 2240 8344 2268 8375
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2406 8344 2412 8356
rect 2240 8316 2412 8344
rect 2406 8304 2412 8316
rect 2464 8344 2470 8356
rect 2884 8344 2912 8452
rect 3513 8449 3525 8452
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 5074 8480 5080 8492
rect 4571 8452 5080 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5184 8480 5212 8511
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 5316 8520 5365 8548
rect 5316 8508 5322 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 5353 8511 5411 8517
rect 5537 8551 5595 8557
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 5644 8548 5672 8576
rect 6380 8548 6408 8576
rect 7006 8548 7012 8560
rect 5583 8520 6408 8548
rect 6748 8520 7012 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 5626 8480 5632 8492
rect 5184 8452 5632 8480
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 6748 8489 6776 8520
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 6135 8452 6745 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 7944 8480 7972 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12434 8616 12440 8628
rect 12115 8588 12440 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 13998 8548 14004 8560
rect 9355 8520 14004 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 13998 8508 14004 8520
rect 14056 8508 14062 8560
rect 6733 8443 6791 8449
rect 6840 8452 7972 8480
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 4062 8412 4068 8424
rect 3743 8384 4068 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 2464 8316 2912 8344
rect 3053 8347 3111 8353
rect 2464 8304 2470 8316
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3237 8347 3295 8353
rect 3237 8344 3249 8347
rect 3099 8316 3249 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3237 8313 3249 8316
rect 3283 8313 3295 8347
rect 3436 8344 3464 8375
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5736 8412 5764 8443
rect 5810 8412 5816 8424
rect 4755 8384 5672 8412
rect 5736 8384 5816 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 3510 8344 3516 8356
rect 3436 8316 3516 8344
rect 3237 8307 3295 8313
rect 3510 8304 3516 8316
rect 3568 8344 3574 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 3568 8316 4813 8344
rect 3568 8304 3574 8316
rect 4801 8313 4813 8316
rect 4847 8313 4859 8347
rect 5644 8344 5672 8384
rect 5810 8372 5816 8384
rect 5868 8412 5874 8424
rect 6840 8412 6868 8452
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9490 8480 9496 8492
rect 9180 8452 9496 8480
rect 9180 8440 9186 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9766 8480 9772 8492
rect 9723 8452 9772 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10318 8480 10324 8492
rect 10091 8452 10324 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 5868 8384 6868 8412
rect 7015 8415 7073 8421
rect 5868 8372 5874 8384
rect 7015 8381 7027 8415
rect 7061 8381 7073 8415
rect 7015 8375 7073 8381
rect 5718 8344 5724 8356
rect 5644 8316 5724 8344
rect 4801 8307 4859 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7024 8344 7052 8375
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9582 8412 9588 8424
rect 9364 8384 9588 8412
rect 9364 8372 9370 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9876 8412 9904 8443
rect 10318 8440 10324 8452
rect 10376 8480 10382 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10376 8452 11161 8480
rect 10376 8440 10382 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 10134 8412 10140 8424
rect 9876 8384 10140 8412
rect 10134 8372 10140 8384
rect 10192 8412 10198 8424
rect 10192 8384 11100 8412
rect 10192 8372 10198 8384
rect 10870 8344 10876 8356
rect 6880 8316 10876 8344
rect 6880 8304 6886 8316
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 3142 8236 3148 8288
rect 3200 8236 3206 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4764 8248 4997 8276
rect 4764 8236 4770 8248
rect 4985 8245 4997 8248
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7190 8276 7196 8288
rect 6963 8248 7196 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9858 8276 9864 8288
rect 8628 8248 9864 8276
rect 8628 8236 8634 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 11072 8285 11100 8384
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 12176 8412 12204 8443
rect 11848 8384 12204 8412
rect 12268 8412 12296 8443
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13538 8480 13544 8492
rect 12943 8452 13544 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12268 8384 12817 8412
rect 11848 8372 11854 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 12912 8276 12940 8443
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 11103 8248 12940 8276
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 1104 8186 13892 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13892 8186
rect 1104 8112 13892 8134
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 5684 8044 8217 8072
rect 5684 8032 5690 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8444 8044 8953 8072
rect 8444 8032 8450 8044
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 9490 8072 9496 8084
rect 8987 8044 9496 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 9674 8032 9680 8084
rect 9732 8032 9738 8084
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 2832 7976 3065 8004
rect 2832 7964 2838 7976
rect 3053 7973 3065 7976
rect 3099 7973 3111 8007
rect 9306 8004 9312 8016
rect 3053 7967 3111 7973
rect 8312 7976 9312 8004
rect 3068 7936 3096 7967
rect 3418 7936 3424 7948
rect 3068 7908 3424 7936
rect 3418 7896 3424 7908
rect 3476 7936 3482 7948
rect 4614 7936 4620 7948
rect 3476 7908 4620 7936
rect 3476 7896 3482 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 1578 7868 1584 7880
rect 1443 7840 1584 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 8312 7877 8340 7976
rect 9306 7964 9312 7976
rect 9364 8004 9370 8016
rect 9364 7976 9674 8004
rect 9364 7964 9370 7976
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 9646 7936 9674 7976
rect 10870 7964 10876 8016
rect 10928 8004 10934 8016
rect 12158 8004 12164 8016
rect 10928 7976 12164 8004
rect 10928 7964 10934 7976
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 9232 7908 9536 7936
rect 9646 7908 11928 7936
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3200 7840 3341 7868
rect 3200 7828 3206 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 1918 7803 1976 7809
rect 1918 7800 1930 7803
rect 1596 7772 1930 7800
rect 1596 7741 1624 7772
rect 1918 7769 1930 7772
rect 1964 7769 1976 7803
rect 8128 7800 8156 7831
rect 8404 7800 8432 7896
rect 9232 7877 9260 7908
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7864 9367 7871
rect 9355 7837 9444 7864
rect 9309 7836 9444 7837
rect 9309 7831 9367 7836
rect 8128 7772 8432 7800
rect 1918 7763 1976 7769
rect 9140 7744 9168 7831
rect 9416 7800 9444 7836
rect 9508 7812 9536 7908
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 11793 7871 11851 7877
rect 11793 7868 11805 7871
rect 11532 7840 11805 7868
rect 9232 7772 9444 7800
rect 9232 7744 9260 7772
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 11532 7809 11560 7840
rect 11793 7837 11805 7840
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 11900 7868 11928 7908
rect 11974 7868 11980 7880
rect 11900 7840 11980 7868
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 9548 7772 9873 7800
rect 9548 7760 9554 7772
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 9861 7763 9919 7769
rect 9953 7803 10011 7809
rect 9953 7769 9965 7803
rect 9999 7800 10011 7803
rect 10321 7803 10379 7809
rect 9999 7772 10180 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 10152 7744 10180 7772
rect 10321 7769 10333 7803
rect 10367 7800 10379 7803
rect 11149 7803 11207 7809
rect 10367 7772 10916 7800
rect 10367 7769 10379 7772
rect 10321 7763 10379 7769
rect 10888 7744 10916 7772
rect 11149 7769 11161 7803
rect 11195 7800 11207 7803
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 11195 7772 11529 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11517 7763 11575 7769
rect 11701 7803 11759 7809
rect 11701 7769 11713 7803
rect 11747 7800 11759 7803
rect 11900 7800 11928 7840
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 11747 7772 11928 7800
rect 11747 7769 11759 7772
rect 11701 7763 11759 7769
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7701 1639 7735
rect 1581 7695 1639 7701
rect 3142 7692 3148 7744
rect 3200 7692 3206 7744
rect 9122 7692 9128 7744
rect 9180 7692 9186 7744
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 10134 7692 10140 7744
rect 10192 7692 10198 7744
rect 10870 7692 10876 7744
rect 10928 7692 10934 7744
rect 11333 7735 11391 7741
rect 11333 7701 11345 7735
rect 11379 7732 11391 7735
rect 11422 7732 11428 7744
rect 11379 7704 11428 7732
rect 11379 7701 11391 7704
rect 11333 7695 11391 7701
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 12066 7692 12072 7744
rect 12124 7692 12130 7744
rect 1104 7642 13892 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 8658 7642
rect 8710 7590 8722 7642
rect 8774 7590 8786 7642
rect 8838 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 13892 7642
rect 1104 7568 13892 7590
rect 3142 7488 3148 7540
rect 3200 7488 3206 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7006 7528 7012 7540
rect 6963 7500 7012 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 2952 7463 3010 7469
rect 2952 7429 2964 7463
rect 2998 7460 3010 7463
rect 3160 7460 3188 7488
rect 2998 7432 3188 7460
rect 5292 7463 5350 7469
rect 2998 7429 3010 7432
rect 2952 7423 3010 7429
rect 5292 7429 5304 7463
rect 5338 7460 5350 7463
rect 5644 7460 5672 7491
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 8478 7528 8484 7540
rect 7944 7500 8484 7528
rect 7650 7460 7656 7472
rect 5338 7432 5672 7460
rect 5828 7432 7656 7460
rect 5338 7429 5350 7432
rect 5292 7423 5350 7429
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 1728 7364 2697 7392
rect 1728 7352 1734 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 1394 7284 1400 7336
rect 1452 7284 1458 7336
rect 5828 7333 5856 7432
rect 7650 7420 7656 7432
rect 7708 7420 7714 7472
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6089 7395 6147 7401
rect 6089 7361 6101 7395
rect 6135 7392 6147 7395
rect 6914 7392 6920 7404
rect 6135 7364 6920 7392
rect 6135 7361 6147 7364
rect 6089 7355 6147 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7944 7401 7972 7500
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9364 7500 9597 7528
rect 9364 7488 9370 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 11238 7488 11244 7540
rect 11296 7488 11302 7540
rect 12158 7488 12164 7540
rect 12216 7488 12222 7540
rect 9122 7460 9128 7472
rect 8312 7432 9128 7460
rect 8312 7401 8340 7432
rect 9122 7420 9128 7432
rect 9180 7460 9186 7472
rect 9180 7432 9904 7460
rect 9180 7420 9186 7432
rect 7469 7395 7527 7401
rect 7469 7361 7481 7395
rect 7515 7392 7527 7395
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7515 7364 7941 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8297 7355 8355 7361
rect 8496 7364 8861 7392
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 5813 7287 5871 7293
rect 5920 7296 6009 7324
rect 1412 7188 1440 7284
rect 3988 7228 4200 7256
rect 3988 7188 4016 7228
rect 1412 7160 4016 7188
rect 4062 7148 4068 7200
rect 4120 7148 4126 7200
rect 4172 7197 4200 7228
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 5920 7188 5948 7296
rect 5997 7293 6009 7296
rect 6043 7293 6055 7327
rect 5997 7287 6055 7293
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 8496 7256 8524 7364
rect 8849 7361 8861 7364
rect 8895 7392 8907 7395
rect 8895 7364 9168 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 7116 7228 8524 7256
rect 7116 7197 7144 7228
rect 4203 7160 5948 7188
rect 7101 7191 7159 7197
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 7101 7157 7113 7191
rect 7147 7157 7159 7191
rect 9140 7188 9168 7364
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9876 7401 9904 7432
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10321 7463 10379 7469
rect 10321 7460 10333 7463
rect 10100 7432 10333 7460
rect 10100 7420 10106 7432
rect 10321 7429 10333 7432
rect 10367 7460 10379 7463
rect 11256 7460 11284 7488
rect 10367 7432 11100 7460
rect 11256 7432 11928 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9272 7364 9413 7392
rect 9272 7352 9278 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10134 7392 10140 7404
rect 9907 7364 10140 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9416 7256 9444 7355
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10192 7364 10517 7392
rect 10192 7352 10198 7364
rect 10505 7361 10517 7364
rect 10551 7392 10563 7395
rect 10686 7392 10692 7404
rect 10551 7364 10692 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9548 7296 9781 7324
rect 9548 7284 9554 7296
rect 9769 7293 9781 7296
rect 9815 7324 9827 7327
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 9815 7296 10793 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 9416 7228 10333 7256
rect 10321 7225 10333 7228
rect 10367 7256 10379 7259
rect 10870 7256 10876 7268
rect 10367 7228 10876 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 10870 7216 10876 7228
rect 10928 7256 10934 7268
rect 10980 7256 11008 7355
rect 10928 7228 11008 7256
rect 10928 7216 10934 7228
rect 11072 7200 11100 7432
rect 11900 7401 11928 7432
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11164 7364 11529 7392
rect 11164 7265 11192 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12032 7364 12081 7392
rect 12032 7352 12038 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 13285 7395 13343 7401
rect 13285 7361 13297 7395
rect 13331 7392 13343 7395
rect 13446 7392 13452 7404
rect 13331 7364 13452 7392
rect 13331 7361 13343 7364
rect 13285 7355 13343 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13538 7284 13544 7336
rect 13596 7284 13602 7336
rect 11149 7259 11207 7265
rect 11149 7225 11161 7259
rect 11195 7225 11207 7259
rect 11149 7219 11207 7225
rect 9582 7188 9588 7200
rect 9140 7160 9588 7188
rect 7101 7151 7159 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11054 7188 11060 7200
rect 11011 7160 11060 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11698 7148 11704 7200
rect 11756 7148 11762 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 12032 7160 12081 7188
rect 12032 7148 12038 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 1104 7098 13892 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13892 7098
rect 1104 7024 13892 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 6822 6984 6828 6996
rect 4120 6956 6828 6984
rect 4120 6944 4126 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7156 6956 7481 6984
rect 7156 6944 7162 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 7469 6947 7527 6953
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 9401 6987 9459 6993
rect 7708 6956 9352 6984
rect 7708 6944 7714 6956
rect 5537 6919 5595 6925
rect 5537 6916 5549 6919
rect 4540 6888 5549 6916
rect 4540 6792 4568 6888
rect 5537 6885 5549 6888
rect 5583 6916 5595 6919
rect 5902 6916 5908 6928
rect 5583 6888 5908 6916
rect 5583 6885 5595 6888
rect 5537 6879 5595 6885
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 7929 6919 7987 6925
rect 7929 6885 7941 6919
rect 7975 6916 7987 6919
rect 9214 6916 9220 6928
rect 7975 6888 9220 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 9324 6916 9352 6956
rect 9401 6953 9413 6987
rect 9447 6984 9459 6987
rect 9582 6984 9588 6996
rect 9447 6956 9588 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 9582 6944 9588 6956
rect 9640 6984 9646 6996
rect 10042 6984 10048 6996
rect 9640 6956 10048 6984
rect 9640 6944 9646 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 11698 6916 11704 6928
rect 9324 6888 11704 6916
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 4939 6820 5396 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5368 6792 5396 6820
rect 5460 6820 6101 6848
rect 5460 6792 5488 6820
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 6089 6811 6147 6817
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 11974 6848 11980 6860
rect 7616 6820 8064 6848
rect 7616 6808 7622 6820
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 5074 6740 5080 6792
rect 5132 6740 5138 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6178 6780 6184 6792
rect 5951 6752 6184 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6356 6783 6414 6789
rect 6356 6749 6368 6783
rect 6402 6780 6414 6783
rect 6914 6780 6920 6792
rect 6402 6752 6920 6780
rect 6402 6749 6414 6752
rect 6356 6743 6414 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 8036 6789 8064 6820
rect 8496 6820 11980 6848
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7156 6752 7757 6780
rect 7156 6740 7162 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 5368 6712 5396 6740
rect 5813 6715 5871 6721
rect 5813 6712 5825 6715
rect 5368 6684 5825 6712
rect 5813 6681 5825 6684
rect 5859 6681 5871 6715
rect 8496 6712 8524 6820
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8588 6752 8953 6780
rect 8588 6724 8616 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9272 6752 9321 6780
rect 9272 6740 9278 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 9539 6752 9573 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 5813 6675 5871 6681
rect 7392 6684 8524 6712
rect 7392 6656 7420 6684
rect 8570 6672 8576 6724
rect 8628 6672 8634 6724
rect 9508 6712 9536 6743
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10704 6789 10732 6820
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10928 6752 10977 6780
rect 10928 6740 10934 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 11112 6752 11161 6780
rect 11112 6740 11118 6752
rect 11149 6749 11161 6752
rect 11195 6780 11207 6783
rect 11195 6752 11836 6780
rect 11195 6749 11207 6752
rect 11149 6743 11207 6749
rect 9048 6684 10732 6712
rect 4246 6604 4252 6656
rect 4304 6604 4310 6656
rect 5258 6604 5264 6656
rect 5316 6604 5322 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 8205 6647 8263 6653
rect 8205 6613 8217 6647
rect 8251 6644 8263 6647
rect 9048 6644 9076 6684
rect 10704 6656 10732 6684
rect 11808 6656 11836 6752
rect 8251 6616 9076 6644
rect 9125 6647 9183 6653
rect 8251 6613 8263 6616
rect 8205 6607 8263 6613
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9398 6644 9404 6656
rect 9171 6616 9404 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10594 6644 10600 6656
rect 9732 6616 10600 6644
rect 9732 6604 9738 6616
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10686 6604 10692 6656
rect 10744 6604 10750 6656
rect 11054 6604 11060 6656
rect 11112 6604 11118 6656
rect 11790 6604 11796 6656
rect 11848 6604 11854 6656
rect 1104 6554 13892 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 8658 6554
rect 8710 6502 8722 6554
rect 8774 6502 8786 6554
rect 8838 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 13892 6554
rect 1104 6480 13892 6502
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4430 6440 4436 6452
rect 4203 6412 4436 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 7745 6443 7803 6449
rect 7745 6440 7757 6443
rect 7616 6412 7757 6440
rect 7616 6400 7622 6412
rect 7745 6409 7757 6412
rect 7791 6409 7803 6443
rect 7745 6403 7803 6409
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9490 6440 9496 6452
rect 9088 6412 9496 6440
rect 9088 6400 9094 6412
rect 9490 6400 9496 6412
rect 9548 6440 9554 6452
rect 9548 6412 10272 6440
rect 9548 6400 9554 6412
rect 4341 6375 4399 6381
rect 4341 6372 4353 6375
rect 2148 6344 4353 6372
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 2148 6313 2176 6344
rect 4341 6341 4353 6344
rect 4387 6372 4399 6375
rect 5442 6372 5448 6384
rect 4387 6344 5448 6372
rect 4387 6341 4399 6344
rect 4341 6335 4399 6341
rect 5442 6332 5448 6344
rect 5500 6372 5506 6384
rect 7834 6372 7840 6384
rect 5500 6344 6408 6372
rect 5500 6332 5506 6344
rect 2406 6313 2412 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1728 6276 2145 6304
rect 1728 6264 1734 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2400 6267 2412 6313
rect 2406 6264 2412 6267
rect 2464 6264 2470 6316
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 3528 6276 3617 6304
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3528 6109 3556 6276
rect 3605 6273 3617 6276
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 3804 6236 3832 6267
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4062 6304 4068 6316
rect 4019 6276 4068 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 6380 6313 6408 6344
rect 6564 6344 7840 6372
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6564 6304 6592 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 9048 6372 9076 6400
rect 8404 6344 9076 6372
rect 6365 6267 6423 6273
rect 6472 6276 6592 6304
rect 6632 6307 6690 6313
rect 4172 6236 4200 6264
rect 3804 6208 4200 6236
rect 6104 6236 6132 6267
rect 6472 6236 6500 6276
rect 6632 6273 6644 6307
rect 6678 6304 6690 6307
rect 7190 6304 7196 6316
rect 6678 6276 7196 6304
rect 6678 6273 6690 6276
rect 6632 6267 6690 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 8404 6313 8432 6344
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9364 6344 10057 6372
rect 9364 6332 9370 6344
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7800 6276 8033 6304
rect 7800 6264 7806 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8662 6304 8668 6316
rect 8619 6276 8668 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 6104 6208 6500 6236
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 3200 6072 3525 6100
rect 3200 6060 3206 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 8220 6100 8248 6267
rect 8662 6264 8668 6276
rect 8720 6304 8726 6316
rect 9214 6304 9220 6316
rect 8720 6276 9220 6304
rect 8720 6264 8726 6276
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 10244 6313 10272 6412
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10652 6412 11192 6440
rect 10652 6400 10658 6412
rect 10336 6344 11008 6372
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 8297 6239 8355 6245
rect 8297 6205 8309 6239
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8312 6168 8340 6199
rect 9582 6168 9588 6180
rect 8312 6140 9588 6168
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 9784 6112 9812 6267
rect 9876 6236 9904 6267
rect 10336 6245 10364 6344
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10686 6304 10692 6316
rect 10459 6276 10692 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10520 6248 10548 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10980 6313 11008 6344
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 11164 6304 11192 6412
rect 11790 6400 11796 6452
rect 11848 6400 11854 6452
rect 11103 6276 11192 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 10321 6239 10379 6245
rect 10321 6236 10333 6239
rect 9876 6208 10333 6236
rect 9876 6112 9904 6208
rect 10321 6205 10333 6208
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 10502 6196 10508 6248
rect 10560 6196 10566 6248
rect 8386 6100 8392 6112
rect 8220 6072 8392 6100
rect 3513 6063 3571 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8536 6072 8769 6100
rect 8536 6060 8542 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9766 6100 9772 6112
rect 9723 6072 9772 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9858 6060 9864 6112
rect 9916 6060 9922 6112
rect 10042 6060 10048 6112
rect 10100 6060 10106 6112
rect 10594 6060 10600 6112
rect 10652 6060 10658 6112
rect 10888 6100 10916 6267
rect 11330 6264 11336 6316
rect 11388 6264 11394 6316
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12906 6307 12964 6313
rect 12906 6304 12918 6307
rect 12492 6276 12918 6304
rect 12492 6264 12498 6276
rect 12906 6273 12918 6276
rect 12952 6273 12964 6307
rect 12906 6267 12964 6273
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 13538 6304 13544 6316
rect 13219 6276 13544 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 11422 6236 11428 6248
rect 11287 6208 11428 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 11054 6100 11060 6112
rect 10888 6072 11060 6100
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 1104 6010 13892 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13892 6010
rect 1104 5936 13892 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2464 5868 2605 5896
rect 2464 5856 2470 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 4893 5899 4951 5905
rect 4893 5865 4905 5899
rect 4939 5896 4951 5899
rect 5074 5896 5080 5908
rect 4939 5868 5080 5896
rect 4939 5865 4951 5868
rect 4893 5859 4951 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5500 5868 6408 5896
rect 5500 5856 5506 5868
rect 4264 5828 4292 5856
rect 2792 5800 4292 5828
rect 2792 5701 2820 5800
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4430 5692 4436 5704
rect 4387 5664 4436 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4614 5652 4620 5704
rect 4672 5652 4678 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4982 5692 4988 5704
rect 4755 5664 4988 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5276 5692 5304 5856
rect 6380 5769 6408 5868
rect 7190 5856 7196 5908
rect 7248 5856 7254 5908
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 8386 5856 8392 5908
rect 8444 5856 8450 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9180 5868 10548 5896
rect 9180 5856 9186 5868
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 8404 5760 8432 5856
rect 10520 5840 10548 5868
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 13538 5896 13544 5908
rect 11756 5868 13544 5896
rect 11756 5856 11762 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 9309 5831 9367 5837
rect 9309 5797 9321 5831
rect 9355 5797 9367 5831
rect 9309 5791 9367 5797
rect 9324 5760 9352 5791
rect 10042 5788 10048 5840
rect 10100 5788 10106 5840
rect 10502 5788 10508 5840
rect 10560 5788 10566 5840
rect 12434 5788 12440 5840
rect 12492 5788 12498 5840
rect 6365 5723 6423 5729
rect 8220 5732 9444 5760
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 5276 5664 6653 5692
rect 6641 5661 6653 5664
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 7742 5692 7748 5704
rect 7699 5664 7748 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 4525 5627 4583 5633
rect 4525 5624 4537 5627
rect 4264 5596 4537 5624
rect 4264 5568 4292 5596
rect 4525 5593 4537 5596
rect 4571 5593 4583 5627
rect 4525 5587 4583 5593
rect 6120 5627 6178 5633
rect 6120 5593 6132 5627
rect 6166 5624 6178 5627
rect 7300 5624 7328 5655
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8220 5701 8248 5732
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8662 5692 8668 5704
rect 8343 5664 8668 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8128 5624 8156 5655
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9030 5692 9036 5704
rect 8987 5664 9036 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9416 5701 9444 5732
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 10060 5760 10088 5788
rect 9640 5732 9996 5760
rect 10060 5732 12480 5760
rect 9640 5720 9646 5732
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9401 5655 9459 5661
rect 9508 5664 9689 5692
rect 6166 5596 6500 5624
rect 7300 5596 8064 5624
rect 8128 5596 8892 5624
rect 6166 5593 6178 5596
rect 6120 5587 6178 5593
rect 4246 5516 4252 5568
rect 4304 5516 4310 5568
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4488 5528 4997 5556
rect 4488 5516 4494 5528
rect 4985 5525 4997 5528
rect 5031 5556 5043 5559
rect 5258 5556 5264 5568
rect 5031 5528 5264 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 6472 5565 6500 5596
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5525 6515 5559
rect 6457 5519 6515 5525
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7607 5528 7941 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 8036 5556 8064 5596
rect 8386 5556 8392 5568
rect 8036 5528 8392 5556
rect 7929 5519 7987 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8864 5556 8892 5596
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 9508 5624 9536 5664
rect 9677 5661 9689 5664
rect 9723 5692 9735 5695
rect 9858 5692 9864 5704
rect 9723 5664 9864 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 9968 5692 9996 5732
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 9968 5664 10333 5692
rect 10321 5661 10333 5664
rect 10367 5661 10379 5695
rect 10321 5655 10379 5661
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 12158 5692 12164 5704
rect 11940 5664 12164 5692
rect 11940 5652 11946 5664
rect 12158 5652 12164 5664
rect 12216 5692 12222 5704
rect 12452 5701 12480 5732
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 12216 5664 12265 5692
rect 12216 5652 12222 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12449 5695 12507 5701
rect 12449 5661 12461 5695
rect 12495 5661 12507 5695
rect 12449 5655 12507 5661
rect 9232 5596 9536 5624
rect 9585 5627 9643 5633
rect 9232 5556 9260 5596
rect 9585 5593 9597 5627
rect 9631 5624 9643 5627
rect 9766 5624 9772 5636
rect 9631 5596 9772 5624
rect 9631 5593 9643 5596
rect 9585 5587 9643 5593
rect 9766 5584 9772 5596
rect 9824 5624 9830 5636
rect 10042 5624 10048 5636
rect 9824 5596 10048 5624
rect 9824 5584 9830 5596
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 8864 5528 9260 5556
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9364 5528 9505 5556
rect 9364 5516 9370 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 11698 5516 11704 5568
rect 11756 5516 11762 5568
rect 1104 5466 13892 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 8658 5466
rect 8710 5414 8722 5466
rect 8774 5414 8786 5466
rect 8838 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 13892 5466
rect 1104 5392 13892 5414
rect 4246 5352 4252 5364
rect 3804 5324 4252 5352
rect 2216 5287 2274 5293
rect 2216 5253 2228 5287
rect 2262 5284 2274 5287
rect 2406 5284 2412 5296
rect 2262 5256 2412 5284
rect 2262 5253 2274 5256
rect 2216 5247 2274 5253
rect 2406 5244 2412 5256
rect 2464 5244 2470 5296
rect 3804 5293 3832 5324
rect 4246 5312 4252 5324
rect 4304 5352 4310 5364
rect 4614 5352 4620 5364
rect 4304 5324 4620 5352
rect 4304 5312 4310 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 10807 5355 10865 5361
rect 9646 5324 10732 5352
rect 3789 5287 3847 5293
rect 3789 5253 3801 5287
rect 3835 5253 3847 5287
rect 5994 5284 6000 5296
rect 3789 5247 3847 5253
rect 3896 5256 6000 5284
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 3896 5225 3924 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 9646 5284 9674 5324
rect 7208 5256 9674 5284
rect 9937 5287 9995 5293
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1728 5188 1961 5216
rect 1728 5176 1734 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 1949 5179 2007 5185
rect 3344 5188 3617 5216
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 3344 5021 3372 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 4062 5216 4068 5228
rect 4019 5188 4068 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4172 5188 4445 5216
rect 4172 5089 4200 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 7208 5225 7236 5256
rect 9937 5253 9949 5287
rect 9983 5284 9995 5287
rect 10137 5287 10195 5293
rect 9983 5256 10088 5284
rect 9983 5253 9995 5256
rect 9937 5247 9995 5253
rect 10060 5228 10088 5256
rect 10137 5253 10149 5287
rect 10183 5284 10195 5287
rect 10502 5284 10508 5296
rect 10183 5256 10364 5284
rect 10183 5253 10195 5256
rect 10137 5247 10195 5253
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7607 5188 9812 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 4580 5120 4629 5148
rect 4580 5108 4586 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 7024 5148 7052 5179
rect 7024 5120 7236 5148
rect 4617 5111 4675 5117
rect 4157 5083 4215 5089
rect 4157 5049 4169 5083
rect 4203 5049 4215 5083
rect 4157 5043 4215 5049
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 6917 5083 6975 5089
rect 6917 5080 6929 5083
rect 6788 5052 6929 5080
rect 6788 5040 6794 5052
rect 6917 5049 6929 5052
rect 6963 5049 6975 5083
rect 6917 5043 6975 5049
rect 7208 5024 7236 5120
rect 9784 5089 9812 5188
rect 10042 5176 10048 5228
rect 10100 5176 10106 5228
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 10336 5157 10364 5256
rect 10428 5256 10508 5284
rect 10428 5225 10456 5256
rect 10502 5244 10508 5256
rect 10560 5284 10566 5296
rect 10597 5287 10655 5293
rect 10597 5284 10609 5287
rect 10560 5256 10609 5284
rect 10560 5244 10566 5256
rect 10597 5253 10609 5256
rect 10643 5253 10655 5287
rect 10704 5284 10732 5324
rect 10807 5321 10819 5355
rect 10853 5352 10865 5355
rect 11054 5352 11060 5364
rect 10853 5324 11060 5352
rect 10853 5321 10865 5324
rect 10807 5315 10865 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11793 5287 11851 5293
rect 10704 5256 11744 5284
rect 10597 5247 10655 5253
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11112 5188 11529 5216
rect 11112 5176 11118 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11609 5219 11667 5225
rect 11609 5185 11621 5219
rect 11655 5185 11667 5219
rect 11609 5179 11667 5185
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9916 5120 10333 5148
rect 9916 5108 9922 5120
rect 10321 5117 10333 5120
rect 10367 5148 10379 5151
rect 11624 5148 11652 5179
rect 10367 5120 11652 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 9769 5083 9827 5089
rect 9769 5049 9781 5083
rect 9815 5049 9827 5083
rect 9769 5043 9827 5049
rect 10244 5052 10824 5080
rect 10244 5024 10272 5052
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 2372 4984 3341 5012
rect 2372 4972 2378 4984
rect 3329 4981 3341 4984
rect 3375 4981 3387 5015
rect 3329 4975 3387 4981
rect 4246 4972 4252 5024
rect 4304 4972 4310 5024
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5537 5015 5595 5021
rect 5537 5012 5549 5015
rect 5500 4984 5549 5012
rect 5500 4972 5506 4984
rect 5537 4981 5549 4984
rect 5583 4981 5595 5015
rect 5537 4975 5595 4981
rect 7190 4972 7196 5024
rect 7248 5012 7254 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7248 4984 7389 5012
rect 7248 4972 7254 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 7377 4975 7435 4981
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10226 5012 10232 5024
rect 9999 4984 10232 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10796 5021 10824 5052
rect 10962 5040 10968 5092
rect 11020 5040 11026 5092
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 4981 10839 5015
rect 11716 5012 11744 5256
rect 11793 5253 11805 5287
rect 11839 5284 11851 5287
rect 13078 5284 13084 5296
rect 11839 5256 13084 5284
rect 11839 5253 11851 5256
rect 11793 5247 11851 5253
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11808 5188 11897 5216
rect 11808 5089 11836 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12066 5216 12072 5228
rect 12023 5188 12072 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 11992 5148 12020 5179
rect 12066 5176 12072 5188
rect 12124 5176 12130 5228
rect 11900 5120 12020 5148
rect 11793 5083 11851 5089
rect 11793 5049 11805 5083
rect 11839 5049 11851 5083
rect 11793 5043 11851 5049
rect 11900 5012 11928 5120
rect 12158 5108 12164 5160
rect 12216 5108 12222 5160
rect 11716 4984 11928 5012
rect 10781 4975 10839 4981
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 12032 4984 12081 5012
rect 12032 4972 12038 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 12069 4975 12127 4981
rect 1104 4922 13892 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13892 4922
rect 1104 4848 13892 4870
rect 2406 4768 2412 4820
rect 2464 4768 2470 4820
rect 4246 4808 4252 4820
rect 2746 4780 4252 4808
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2746 4604 2774 4780
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 8297 4811 8355 4817
rect 7892 4780 8156 4808
rect 7892 4768 7898 4780
rect 8128 4681 8156 4780
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8478 4808 8484 4820
rect 8343 4780 8484 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9640 4780 9965 4808
rect 9640 4768 9646 4780
rect 9953 4777 9965 4780
rect 9999 4808 10011 4811
rect 9999 4780 10180 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 8570 4700 8576 4752
rect 8628 4740 8634 4752
rect 9309 4743 9367 4749
rect 9309 4740 9321 4743
rect 8628 4712 9321 4740
rect 8628 4700 8634 4712
rect 9309 4709 9321 4712
rect 9355 4740 9367 4743
rect 9493 4743 9551 4749
rect 9493 4740 9505 4743
rect 9355 4712 9505 4740
rect 9355 4709 9367 4712
rect 9309 4703 9367 4709
rect 9493 4709 9505 4712
rect 9539 4709 9551 4743
rect 9858 4740 9864 4752
rect 9493 4703 9551 4709
rect 9784 4712 9864 4740
rect 8113 4675 8171 4681
rect 3804 4644 4844 4672
rect 3804 4616 3832 4644
rect 2639 4576 2774 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4816 4613 4844 4644
rect 8113 4641 8125 4675
rect 8159 4641 8171 4675
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8113 4635 8171 4641
rect 8404 4644 8953 4672
rect 8404 4616 8432 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 9674 4672 9680 4684
rect 8941 4635 8999 4641
rect 9140 4644 9680 4672
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 4982 4604 4988 4616
rect 4939 4576 4988 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 4540 4468 4568 4567
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5166 4564 5172 4616
rect 5224 4564 5230 4616
rect 5442 4613 5448 4616
rect 5436 4604 5448 4613
rect 5403 4576 5448 4604
rect 5436 4567 5448 4576
rect 5442 4564 5448 4567
rect 5500 4564 5506 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7432 4576 8033 4604
rect 7432 4564 7438 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 9140 4613 9168 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9784 4681 9812 4712
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4641 9827 4675
rect 9769 4635 9827 4641
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 4614 4496 4620 4548
rect 4672 4536 4678 4548
rect 4709 4539 4767 4545
rect 4709 4536 4721 4539
rect 4672 4508 4721 4536
rect 4672 4496 4678 4508
rect 4709 4505 4721 4508
rect 4755 4505 4767 4539
rect 7098 4536 7104 4548
rect 4709 4499 4767 4505
rect 4816 4508 7104 4536
rect 4816 4468 4844 4508
rect 4540 4440 4844 4468
rect 5074 4428 5080 4480
rect 5132 4428 5138 4480
rect 6564 4477 6592 4508
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 7776 4539 7834 4545
rect 7776 4505 7788 4539
rect 7822 4536 7834 4539
rect 7926 4536 7932 4548
rect 7822 4508 7932 4536
rect 7822 4505 7834 4508
rect 7776 4499 7834 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8662 4536 8668 4548
rect 8036 4508 8668 4536
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 6641 4471 6699 4477
rect 6641 4437 6653 4471
rect 6687 4468 6699 4471
rect 8036 4468 8064 4508
rect 8662 4496 8668 4508
rect 8720 4536 8726 4548
rect 8772 4536 8800 4567
rect 9398 4564 9404 4616
rect 9456 4564 9462 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10152 4604 10180 4780
rect 13078 4768 13084 4820
rect 13136 4768 13142 4820
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10652 4644 10977 4672
rect 10652 4632 10658 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 10873 4607 10931 4613
rect 10873 4604 10885 4607
rect 10152 4576 10885 4604
rect 8720 4508 8800 4536
rect 8720 4496 8726 4508
rect 6687 4440 8064 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 8110 4428 8116 4480
rect 8168 4428 8174 4480
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 10152 4468 10180 4576
rect 10873 4573 10885 4576
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11698 4604 11704 4616
rect 11112 4576 11704 4604
rect 11112 4564 11118 4576
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11974 4613 11980 4616
rect 11968 4604 11980 4613
rect 11935 4576 11980 4604
rect 11968 4567 11980 4576
rect 11974 4564 11980 4567
rect 12032 4564 12038 4616
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 11514 4536 11520 4548
rect 10827 4508 11520 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 8619 4440 10180 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 1104 4378 13892 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 8658 4378
rect 8710 4326 8722 4378
rect 8774 4326 8786 4378
rect 8838 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 13892 4378
rect 1104 4304 13892 4326
rect 4614 4264 4620 4276
rect 3988 4236 4620 4264
rect 3988 4196 4016 4236
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 5074 4224 5080 4276
rect 5132 4224 5138 4276
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 5718 4264 5724 4276
rect 5675 4236 5724 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 8110 4224 8116 4276
rect 8168 4224 8174 4276
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8386 4264 8392 4276
rect 8343 4236 8392 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8478 4224 8484 4276
rect 8536 4224 8542 4276
rect 10410 4224 10416 4276
rect 10468 4224 10474 4276
rect 3896 4168 4016 4196
rect 4080 4168 5028 4196
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 2406 4137 2412 4140
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 1728 4100 2145 4128
rect 1728 4088 1734 4100
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2400 4091 2412 4137
rect 2406 4088 2412 4091
rect 2464 4088 2470 4140
rect 3896 4137 3924 4168
rect 4080 4140 4108 4168
rect 5000 4140 5028 4168
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3620 4100 3709 4128
rect 3620 3936 3648 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4062 4088 4068 4140
rect 4120 4088 4126 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4264 4100 4537 4128
rect 4264 4001 4292 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5092 4128 5120 4224
rect 7834 4196 7840 4208
rect 5552 4168 7840 4196
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5092 4100 5457 4128
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5350 4060 5356 4072
rect 5307 4032 5356 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 4249 3995 4307 4001
rect 4249 3961 4261 3995
rect 4295 3961 4307 3995
rect 4249 3955 4307 3961
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 4724 3992 4752 4023
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5552 4060 5580 4168
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 5460 4032 5580 4060
rect 7852 4060 7880 4156
rect 8128 4137 8156 4224
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8496 4128 8524 4224
rect 10428 4196 10456 4224
rect 10244 4168 10456 4196
rect 10244 4137 10272 4168
rect 8435 4100 8524 4128
rect 10229 4131 10287 4137
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10459 4100 10609 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 7852 4032 10057 4060
rect 5460 3992 5488 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 4580 3964 5488 3992
rect 4580 3952 4586 3964
rect 7926 3952 7932 4004
rect 7984 3992 7990 4004
rect 8113 3995 8171 4001
rect 8113 3992 8125 3995
rect 7984 3964 8125 3992
rect 7984 3952 7990 3964
rect 8113 3961 8125 3964
rect 8159 3961 8171 3995
rect 8113 3955 8171 3961
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 12158 3992 12164 4004
rect 8444 3964 12164 3992
rect 8444 3952 8450 3964
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 3513 3927 3571 3933
rect 3513 3893 3525 3927
rect 3559 3924 3571 3927
rect 3602 3924 3608 3936
rect 3559 3896 3608 3924
rect 3559 3893 3571 3896
rect 3513 3887 3571 3893
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 10778 3884 10784 3936
rect 10836 3884 10842 3936
rect 1104 3834 13892 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13892 3834
rect 1104 3760 13892 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 2501 3723 2559 3729
rect 2501 3720 2513 3723
rect 2464 3692 2513 3720
rect 2464 3680 2470 3692
rect 2501 3689 2513 3692
rect 2547 3689 2559 3723
rect 4338 3720 4344 3732
rect 2501 3683 2559 3689
rect 2700 3692 4344 3720
rect 2700 3525 2728 3692
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 11572 3692 11989 3720
rect 11572 3680 11578 3692
rect 11977 3689 11989 3692
rect 12023 3689 12035 3723
rect 11977 3683 12035 3689
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 13504 3692 13553 3720
rect 13504 3680 13510 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 13541 3683 13599 3689
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 9122 3652 9128 3664
rect 8527 3624 9128 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 3292 3556 5120 3584
rect 3292 3544 3298 3556
rect 4062 3525 4068 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 4041 3519 4068 3525
rect 4041 3485 4053 3519
rect 4041 3479 4068 3485
rect 4062 3476 4068 3479
rect 4120 3476 4126 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4172 3448 4200 3479
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5092 3525 5120 3556
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5224 3556 6101 3584
rect 5224 3544 5230 3556
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 7432 3556 10609 3584
rect 7432 3544 7438 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5994 3516 6000 3528
rect 5399 3488 6000 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 6972 3488 7573 3516
rect 6972 3476 6978 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7742 3476 7748 3528
rect 7800 3476 7806 3528
rect 7834 3476 7840 3528
rect 7892 3476 7898 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8711 3488 8953 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 3752 3420 4200 3448
rect 4249 3451 4307 3457
rect 3752 3408 3758 3420
rect 4249 3417 4261 3451
rect 4295 3448 4307 3451
rect 4614 3448 4620 3460
rect 4295 3420 4620 3448
rect 4295 3417 4307 3420
rect 4249 3411 4307 3417
rect 4614 3408 4620 3420
rect 4672 3448 4678 3460
rect 5169 3451 5227 3457
rect 5169 3448 5181 3451
rect 4672 3420 5181 3448
rect 4672 3408 4678 3420
rect 5169 3417 5181 3420
rect 5215 3417 5227 3451
rect 5169 3411 5227 3417
rect 6356 3451 6414 3457
rect 6356 3417 6368 3451
rect 6402 3448 6414 3451
rect 6638 3448 6644 3460
rect 6402 3420 6644 3448
rect 6402 3417 6414 3420
rect 6356 3411 6414 3417
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 4798 3340 4804 3392
rect 4856 3340 4862 3392
rect 5184 3380 5212 3411
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 6730 3408 6736 3460
rect 6788 3408 6794 3460
rect 8294 3408 8300 3460
rect 8352 3408 8358 3460
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 8757 3451 8815 3457
rect 8757 3448 8769 3451
rect 8628 3420 8769 3448
rect 8628 3408 8634 3420
rect 8757 3417 8769 3420
rect 8803 3417 8815 3451
rect 8956 3448 8984 3479
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9263 3488 9628 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 8956 3420 9321 3448
rect 8757 3411 8815 3417
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 6748 3380 6776 3408
rect 9600 3392 9628 3488
rect 5184 3352 6776 3380
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 7064 3352 7481 3380
rect 7064 3340 7070 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 9582 3340 9588 3392
rect 9640 3340 9646 3392
rect 10612 3380 10640 3547
rect 10864 3519 10922 3525
rect 10864 3485 10876 3519
rect 10910 3485 10922 3519
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 10864 3479 10922 3485
rect 11072 3488 12173 3516
rect 10778 3408 10784 3460
rect 10836 3448 10842 3460
rect 10888 3448 10916 3479
rect 10836 3420 10916 3448
rect 10836 3408 10842 3420
rect 11072 3392 11100 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12428 3451 12486 3457
rect 12428 3417 12440 3451
rect 12474 3448 12486 3451
rect 13354 3448 13360 3460
rect 12474 3420 13360 3448
rect 12474 3417 12486 3420
rect 12428 3411 12486 3417
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 11054 3380 11060 3392
rect 10612 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 1104 3290 13892 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 8658 3290
rect 8710 3238 8722 3290
rect 8774 3238 8786 3290
rect 8838 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 13892 3290
rect 1104 3216 13892 3238
rect 4982 3136 4988 3188
rect 5040 3176 5046 3188
rect 5040 3148 5304 3176
rect 5040 3136 5046 3148
rect 5276 3108 5304 3148
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 7742 3176 7748 3188
rect 7147 3148 7748 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 9416 3148 9689 3176
rect 2792 3080 5212 3108
rect 5276 3080 6675 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 2792 3049 2820 3080
rect 3050 3049 3056 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 1728 3012 2789 3040
rect 1728 3000 1734 3012
rect 2777 3009 2789 3012
rect 2823 3040 2835 3043
rect 2823 3012 2877 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 3044 3003 3056 3049
rect 3050 3000 3056 3003
rect 3108 3000 3114 3052
rect 4338 3000 4344 3052
rect 4396 3000 4402 3052
rect 4632 3049 4660 3080
rect 5184 3052 5212 3080
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4873 3043 4931 3049
rect 4873 3040 4885 3043
rect 4617 3003 4675 3009
rect 4724 3012 4885 3040
rect 4724 2972 4752 3012
rect 4873 3009 4885 3012
rect 4919 3009 4931 3043
rect 4873 3003 4931 3009
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6647 3040 6675 3080
rect 6730 3068 6736 3120
rect 6788 3068 6794 3120
rect 6822 3068 6828 3120
rect 6880 3068 6886 3120
rect 7190 3108 7196 3120
rect 6932 3080 7196 3108
rect 6932 3049 6960 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 7644 3111 7702 3117
rect 7644 3077 7656 3111
rect 7690 3108 7702 3111
rect 8312 3108 8340 3136
rect 7690 3080 8340 3108
rect 7690 3077 7702 3080
rect 7644 3071 7702 3077
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6647 3012 6929 3040
rect 6549 3003 6607 3009
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 4540 2944 4752 2972
rect 6564 2972 6592 3003
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7984 3012 8861 3040
rect 7984 3000 7990 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9140 3040 9168 3136
rect 9416 3052 9444 3148
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 9140 3012 9229 3040
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 9398 3000 9404 3052
rect 9456 3000 9462 3052
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3040 9643 3043
rect 10790 3043 10848 3049
rect 10790 3040 10802 3043
rect 9631 3012 10802 3040
rect 9631 3009 9643 3012
rect 9585 3003 9643 3009
rect 10790 3009 10802 3012
rect 10836 3009 10848 3043
rect 10790 3003 10848 3009
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 7024 2972 7052 3000
rect 6564 2944 7052 2972
rect 9125 2975 9183 2981
rect 4540 2913 4568 2944
rect 9125 2941 9137 2975
rect 9171 2972 9183 2975
rect 9306 2972 9312 2984
rect 9171 2944 9312 2972
rect 9171 2941 9183 2944
rect 9125 2935 9183 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 4525 2907 4583 2913
rect 4525 2873 4537 2907
rect 4571 2873 4583 2907
rect 4525 2867 4583 2873
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4430 2836 4436 2848
rect 4203 2808 4436 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 9398 2836 9404 2848
rect 8803 2808 9404 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 9398 2796 9404 2808
rect 9456 2836 9462 2848
rect 9582 2836 9588 2848
rect 9456 2808 9588 2836
rect 9456 2796 9462 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 1104 2746 13892 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13892 2746
rect 1104 2672 13892 2694
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 3108 2604 3157 2632
rect 3108 2592 3114 2604
rect 3145 2601 3157 2604
rect 3191 2601 3203 2635
rect 3145 2595 3203 2601
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4396 2604 4997 2632
rect 4396 2592 4402 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 6638 2592 6644 2644
rect 6696 2592 6702 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7156 2604 8432 2632
rect 7156 2592 7162 2604
rect 5258 2524 5264 2576
rect 5316 2564 5322 2576
rect 8404 2564 8432 2604
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 13354 2592 13360 2644
rect 13412 2592 13418 2644
rect 5316 2536 8340 2564
rect 8404 2536 9628 2564
rect 5316 2524 5322 2536
rect 3142 2496 3148 2508
rect 1596 2468 3148 2496
rect 1596 2437 1624 2468
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3344 2468 3801 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 2314 2388 2320 2440
rect 2372 2388 2378 2440
rect 3344 2437 3372 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4522 2496 4528 2508
rect 4203 2468 4528 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4522 2456 4528 2468
rect 4580 2496 4586 2508
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 4580 2468 5365 2496
rect 4580 2456 4586 2468
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 6914 2496 6920 2508
rect 5353 2459 5411 2465
rect 6840 2468 6920 2496
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3602 2388 3608 2440
rect 3660 2388 3666 2440
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4488 2400 4721 2428
rect 4488 2388 4494 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4856 2400 5181 2428
rect 4856 2388 4862 2400
rect 5169 2397 5181 2400
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 5994 2428 6000 2440
rect 5951 2400 6000 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6840 2437 6868 2468
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7006 2456 7012 2508
rect 7064 2456 7070 2508
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 7024 2428 7052 2456
rect 8312 2437 8340 2536
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 7024 2400 7113 2428
rect 6825 2391 6883 2397
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8628 2400 9045 2428
rect 8628 2388 8634 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9398 2428 9404 2440
rect 9355 2400 9404 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 9600 2437 9628 2536
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9916 2400 10149 2428
rect 9916 2388 9922 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10137 2391 10195 2397
rect 10336 2400 10701 2428
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2360 9275 2363
rect 9508 2360 9536 2388
rect 9263 2332 9536 2360
rect 9263 2329 9275 2332
rect 9217 2323 9275 2329
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 900 2264 1409 2292
rect 900 2252 906 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 2130 2252 2136 2304
rect 2188 2252 2194 2304
rect 3418 2252 3424 2304
rect 3476 2252 3482 2304
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 5718 2252 5724 2304
rect 5776 2252 5782 2304
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6880 2264 6929 2292
rect 6880 2252 6886 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 6917 2255 6975 2261
rect 8110 2252 8116 2304
rect 8168 2252 8174 2304
rect 9398 2252 9404 2304
rect 9456 2252 9462 2304
rect 10336 2301 10364 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11572 2400 11897 2428
rect 11572 2388 11578 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 13078 2388 13084 2440
rect 13136 2388 13142 2440
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 13998 2428 14004 2440
rect 13587 2400 14004 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 10321 2295 10379 2301
rect 10321 2261 10333 2295
rect 10367 2261 10379 2295
rect 10321 2255 10379 2261
rect 10502 2252 10508 2304
rect 10560 2252 10566 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 12894 2252 12900 2304
rect 12952 2252 12958 2304
rect 1104 2202 13892 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 8658 2202
rect 8710 2150 8722 2202
rect 8774 2150 8786 2202
rect 8838 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 13892 2202
rect 1104 2128 13892 2150
<< via1 >>
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 848 14560 900 14612
rect 1768 14560 1820 14612
rect 2872 14560 2924 14612
rect 3884 14560 3936 14612
rect 4896 14560 4948 14612
rect 5908 14560 5960 14612
rect 6920 14560 6972 14612
rect 7840 14560 7892 14612
rect 8944 14560 8996 14612
rect 4712 14424 4764 14476
rect 1768 14356 1820 14408
rect 3056 14356 3108 14408
rect 3516 14356 3568 14408
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 3240 14288 3292 14340
rect 3700 14288 3752 14340
rect 5632 14356 5684 14408
rect 7288 14356 7340 14408
rect 10968 14356 11020 14408
rect 11980 14356 12032 14408
rect 12992 14356 13044 14408
rect 6184 14220 6236 14272
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 12992 14220 13044 14272
rect 2658 14118 2710 14170
rect 2722 14118 2774 14170
rect 2786 14118 2838 14170
rect 2850 14118 2902 14170
rect 2914 14118 2966 14170
rect 2978 14118 3030 14170
rect 8658 14118 8710 14170
rect 8722 14118 8774 14170
rect 8786 14118 8838 14170
rect 8850 14118 8902 14170
rect 8914 14118 8966 14170
rect 8978 14118 9030 14170
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 1584 13948 1636 14000
rect 1400 13880 1452 13932
rect 2412 13880 2464 13932
rect 3424 13880 3476 13932
rect 5540 13948 5592 14000
rect 4896 13880 4948 13932
rect 7472 13880 7524 13932
rect 9496 13923 9548 13932
rect 9496 13889 9514 13923
rect 9514 13889 9548 13923
rect 9496 13880 9548 13889
rect 10416 13880 10468 13932
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 1676 13676 1728 13728
rect 4620 13676 4672 13728
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 7840 13676 7892 13728
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 9404 13676 9456 13728
rect 11796 13744 11848 13796
rect 11152 13676 11204 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 3976 13472 4028 13524
rect 5632 13472 5684 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 7472 13472 7524 13524
rect 4896 13404 4948 13456
rect 1492 13268 1544 13320
rect 1676 13311 1728 13320
rect 1676 13277 1710 13311
rect 1710 13277 1728 13311
rect 1676 13268 1728 13277
rect 3608 13268 3660 13320
rect 5540 13336 5592 13388
rect 7840 13336 7892 13388
rect 4528 13268 4580 13320
rect 4988 13268 5040 13320
rect 5448 13268 5500 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 3332 13132 3384 13184
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 5356 13200 5408 13252
rect 5908 13132 5960 13184
rect 9772 13404 9824 13456
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 8484 13132 8536 13184
rect 10048 13268 10100 13320
rect 10416 13472 10468 13524
rect 10232 13404 10284 13456
rect 11612 13404 11664 13456
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10232 13132 10284 13184
rect 11060 13268 11112 13320
rect 11336 13200 11388 13252
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 11152 13132 11204 13184
rect 11612 13132 11664 13184
rect 11704 13132 11756 13184
rect 11980 13132 12032 13184
rect 2658 13030 2710 13082
rect 2722 13030 2774 13082
rect 2786 13030 2838 13082
rect 2850 13030 2902 13082
rect 2914 13030 2966 13082
rect 2978 13030 3030 13082
rect 8658 13030 8710 13082
rect 8722 13030 8774 13082
rect 8786 13030 8838 13082
rect 8850 13030 8902 13082
rect 8914 13030 8966 13082
rect 8978 13030 9030 13082
rect 3056 12928 3108 12980
rect 3424 12971 3476 12980
rect 3424 12937 3433 12971
rect 3433 12937 3467 12971
rect 3467 12937 3476 12971
rect 3424 12928 3476 12937
rect 3608 12928 3660 12980
rect 4528 12928 4580 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 5908 12928 5960 12980
rect 7380 12928 7432 12980
rect 8024 12928 8076 12980
rect 9772 12928 9824 12980
rect 10692 12928 10744 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 1584 12792 1636 12844
rect 1768 12835 1820 12844
rect 1768 12801 1802 12835
rect 1802 12801 1820 12835
rect 1768 12792 1820 12801
rect 3332 12860 3384 12912
rect 3884 12903 3936 12912
rect 3884 12869 3893 12903
rect 3893 12869 3927 12903
rect 3927 12869 3936 12903
rect 3884 12860 3936 12869
rect 4804 12903 4856 12912
rect 4804 12869 4813 12903
rect 4813 12869 4847 12903
rect 4847 12869 4856 12903
rect 4804 12860 4856 12869
rect 6184 12903 6236 12912
rect 6184 12869 6193 12903
rect 6193 12869 6227 12903
rect 6227 12869 6236 12903
rect 6184 12860 6236 12869
rect 7288 12860 7340 12912
rect 3148 12656 3200 12708
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 4712 12792 4764 12844
rect 5080 12792 5132 12844
rect 4988 12724 5040 12776
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 5448 12724 5500 12776
rect 5724 12724 5776 12776
rect 5816 12656 5868 12708
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 9220 12792 9272 12844
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 11612 12860 11664 12912
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 9588 12724 9640 12776
rect 10600 12835 10652 12844
rect 10600 12801 10614 12835
rect 10614 12801 10648 12835
rect 10648 12801 10652 12835
rect 10600 12792 10652 12801
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 10876 12724 10928 12776
rect 11796 12792 11848 12844
rect 9772 12656 9824 12708
rect 10232 12656 10284 12708
rect 10416 12656 10468 12708
rect 10692 12656 10744 12708
rect 11336 12656 11388 12708
rect 10048 12588 10100 12640
rect 10324 12588 10376 12640
rect 12164 12656 12216 12708
rect 11980 12588 12032 12640
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 1768 12384 1820 12436
rect 2412 12384 2464 12436
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 3056 12316 3108 12368
rect 3240 12316 3292 12368
rect 4712 12316 4764 12368
rect 5356 12316 5408 12368
rect 8668 12384 8720 12436
rect 10784 12384 10836 12436
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 11520 12384 11572 12436
rect 1768 12180 1820 12232
rect 2504 12180 2556 12232
rect 3056 12180 3108 12232
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 9312 12316 9364 12368
rect 4528 12112 4580 12164
rect 6276 12112 6328 12164
rect 8300 12180 8352 12232
rect 8392 12180 8444 12232
rect 9404 12248 9456 12300
rect 9864 12248 9916 12300
rect 9680 12180 9732 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 8484 12112 8536 12164
rect 9505 12155 9557 12164
rect 9505 12121 9539 12155
rect 9539 12121 9557 12155
rect 9505 12112 9557 12121
rect 9772 12112 9824 12164
rect 11060 12180 11112 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 4896 12044 4948 12096
rect 5448 12044 5500 12096
rect 7104 12044 7156 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7840 12044 7892 12096
rect 10600 12112 10652 12164
rect 10416 12044 10468 12096
rect 11152 12044 11204 12096
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 11888 12112 11940 12164
rect 11612 12044 11664 12096
rect 12348 12155 12400 12164
rect 12348 12121 12382 12155
rect 12382 12121 12400 12155
rect 12348 12112 12400 12121
rect 12532 12112 12584 12164
rect 12440 12044 12492 12096
rect 12900 12044 12952 12096
rect 2658 11942 2710 11994
rect 2722 11942 2774 11994
rect 2786 11942 2838 11994
rect 2850 11942 2902 11994
rect 2914 11942 2966 11994
rect 2978 11942 3030 11994
rect 8658 11942 8710 11994
rect 8722 11942 8774 11994
rect 8786 11942 8838 11994
rect 8850 11942 8902 11994
rect 8914 11942 8966 11994
rect 8978 11942 9030 11994
rect 2688 11772 2740 11824
rect 3056 11840 3108 11892
rect 3516 11840 3568 11892
rect 4804 11840 4856 11892
rect 5172 11840 5224 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 5816 11840 5868 11892
rect 8484 11840 8536 11892
rect 9496 11883 9548 11892
rect 1584 11636 1636 11688
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3240 11772 3292 11824
rect 5632 11772 5684 11824
rect 6276 11772 6328 11824
rect 9128 11815 9180 11824
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 2320 11636 2372 11645
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 2964 11636 3016 11688
rect 3792 11704 3844 11756
rect 3148 11568 3200 11620
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6552 11679 6604 11688
rect 6552 11645 6570 11679
rect 6570 11645 6604 11679
rect 6552 11636 6604 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 9128 11781 9137 11815
rect 9137 11781 9171 11815
rect 9171 11781 9180 11815
rect 9128 11772 9180 11781
rect 8392 11704 8444 11756
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 10140 11840 10192 11892
rect 10876 11840 10928 11892
rect 11336 11840 11388 11892
rect 9680 11772 9732 11824
rect 11152 11772 11204 11824
rect 12348 11840 12400 11892
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 10232 11704 10284 11756
rect 10508 11747 10560 11756
rect 8300 11636 8352 11688
rect 9128 11568 9180 11620
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 11060 11704 11112 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 12440 11772 12492 11824
rect 12900 11747 12952 11756
rect 3516 11500 3568 11552
rect 4160 11500 4212 11552
rect 4804 11500 4856 11552
rect 6184 11500 6236 11552
rect 10416 11500 10468 11552
rect 11152 11568 11204 11620
rect 11244 11568 11296 11620
rect 12164 11636 12216 11688
rect 12440 11636 12492 11688
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 11704 11500 11756 11552
rect 12992 11568 13044 11620
rect 12164 11500 12216 11552
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 1676 11296 1728 11348
rect 1768 11296 1820 11348
rect 2412 11296 2464 11348
rect 2504 11296 2556 11348
rect 3056 11296 3108 11348
rect 3240 11296 3292 11348
rect 3700 11296 3752 11348
rect 5080 11296 5132 11348
rect 5632 11296 5684 11348
rect 2688 11228 2740 11280
rect 3332 11228 3384 11280
rect 3516 11228 3568 11280
rect 6368 11296 6420 11348
rect 6736 11296 6788 11348
rect 7380 11296 7432 11348
rect 7840 11296 7892 11348
rect 9128 11296 9180 11348
rect 12164 11296 12216 11348
rect 1768 11092 1820 11144
rect 8116 11228 8168 11280
rect 9496 11228 9548 11280
rect 10508 11228 10560 11280
rect 4160 11092 4212 11144
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 3608 11024 3660 11076
rect 4068 11024 4120 11076
rect 4988 11024 5040 11076
rect 5724 11092 5776 11144
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6184 11092 6236 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 6644 11024 6696 11076
rect 7196 11092 7248 11144
rect 7564 11092 7616 11144
rect 9128 11160 9180 11212
rect 8484 11092 8536 11144
rect 10232 11160 10284 11212
rect 9772 11092 9824 11144
rect 10508 11092 10560 11144
rect 9680 11024 9732 11076
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11244 11092 11296 11144
rect 2964 10956 3016 11008
rect 4620 10999 4672 11008
rect 4620 10965 4629 10999
rect 4629 10965 4663 10999
rect 4663 10965 4672 10999
rect 4620 10956 4672 10965
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 8116 10956 8168 11008
rect 11152 11024 11204 11076
rect 11520 11024 11572 11076
rect 10692 10956 10744 11008
rect 11796 10956 11848 11008
rect 2658 10854 2710 10906
rect 2722 10854 2774 10906
rect 2786 10854 2838 10906
rect 2850 10854 2902 10906
rect 2914 10854 2966 10906
rect 2978 10854 3030 10906
rect 8658 10854 8710 10906
rect 8722 10854 8774 10906
rect 8786 10854 8838 10906
rect 8850 10854 8902 10906
rect 8914 10854 8966 10906
rect 8978 10854 9030 10906
rect 1400 10752 1452 10804
rect 3148 10752 3200 10804
rect 7012 10752 7064 10804
rect 7840 10752 7892 10804
rect 7932 10752 7984 10804
rect 8116 10752 8168 10804
rect 8484 10752 8536 10804
rect 9220 10752 9272 10804
rect 3056 10727 3108 10736
rect 3056 10693 3083 10727
rect 3083 10693 3108 10727
rect 3056 10684 3108 10693
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2780 10616 2832 10668
rect 4068 10684 4120 10736
rect 6736 10616 6788 10668
rect 1492 10591 1544 10600
rect 1492 10557 1501 10591
rect 1501 10557 1535 10591
rect 1535 10557 1544 10591
rect 1492 10548 1544 10557
rect 3700 10548 3752 10600
rect 3976 10548 4028 10600
rect 7564 10548 7616 10600
rect 7748 10616 7800 10668
rect 8392 10548 8444 10600
rect 3608 10480 3660 10532
rect 7748 10480 7800 10532
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 10324 10752 10376 10804
rect 10508 10752 10560 10804
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10048 10548 10100 10600
rect 9404 10523 9456 10532
rect 9404 10489 9413 10523
rect 9413 10489 9447 10523
rect 9447 10489 9456 10523
rect 9404 10480 9456 10489
rect 9588 10480 9640 10532
rect 11060 10752 11112 10804
rect 11980 10752 12032 10804
rect 12532 10752 12584 10804
rect 11244 10684 11296 10736
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 10600 10548 10652 10600
rect 10692 10548 10744 10600
rect 11520 10548 11572 10600
rect 2320 10412 2372 10464
rect 4620 10412 4672 10464
rect 4712 10412 4764 10464
rect 5540 10412 5592 10464
rect 6920 10412 6972 10464
rect 10140 10412 10192 10464
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12808 10412 12860 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 1492 10208 1544 10260
rect 2320 10208 2372 10260
rect 3056 10208 3108 10260
rect 4160 10208 4212 10260
rect 5724 10208 5776 10260
rect 5816 10208 5868 10260
rect 6184 10208 6236 10260
rect 6368 10208 6420 10260
rect 6460 10208 6512 10260
rect 1492 10072 1544 10124
rect 1768 10072 1820 10124
rect 4252 10140 4304 10192
rect 4620 10140 4672 10192
rect 5264 10140 5316 10192
rect 2504 10004 2556 10056
rect 2412 9936 2464 9988
rect 6368 10072 6420 10124
rect 7288 10208 7340 10260
rect 7656 10208 7708 10260
rect 9404 10208 9456 10260
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 10600 10208 10652 10260
rect 11612 10208 11664 10260
rect 11704 10208 11756 10260
rect 12164 10208 12216 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 8944 10140 8996 10192
rect 7472 10072 7524 10124
rect 8484 10072 8536 10124
rect 10048 10140 10100 10192
rect 13544 10140 13596 10192
rect 3608 9936 3660 9988
rect 5080 9936 5132 9988
rect 5816 10004 5868 10056
rect 5448 9936 5500 9988
rect 6092 10004 6144 10056
rect 6644 10004 6696 10056
rect 2780 9868 2832 9920
rect 4528 9868 4580 9920
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 4712 9868 4764 9920
rect 4896 9868 4948 9920
rect 5356 9868 5408 9920
rect 9496 10004 9548 10056
rect 9588 10004 9640 10056
rect 9864 10004 9916 10056
rect 10232 10004 10284 10056
rect 11336 10004 11388 10056
rect 12256 10004 12308 10056
rect 7380 9936 7432 9988
rect 7656 9936 7708 9988
rect 7840 9936 7892 9988
rect 10416 9979 10468 9988
rect 10416 9945 10425 9979
rect 10425 9945 10459 9979
rect 10459 9945 10468 9979
rect 10416 9936 10468 9945
rect 11244 9936 11296 9988
rect 7564 9868 7616 9920
rect 11428 9868 11480 9920
rect 11612 9868 11664 9920
rect 12532 9936 12584 9988
rect 2658 9766 2710 9818
rect 2722 9766 2774 9818
rect 2786 9766 2838 9818
rect 2850 9766 2902 9818
rect 2914 9766 2966 9818
rect 2978 9766 3030 9818
rect 8658 9766 8710 9818
rect 8722 9766 8774 9818
rect 8786 9766 8838 9818
rect 8850 9766 8902 9818
rect 8914 9766 8966 9818
rect 8978 9766 9030 9818
rect 4528 9664 4580 9716
rect 4620 9664 4672 9716
rect 5172 9664 5224 9716
rect 5264 9664 5316 9716
rect 6368 9664 6420 9716
rect 4988 9639 5040 9648
rect 4988 9605 4997 9639
rect 4997 9605 5031 9639
rect 5031 9605 5040 9639
rect 4988 9596 5040 9605
rect 1768 9460 1820 9512
rect 4896 9460 4948 9512
rect 9496 9707 9548 9716
rect 9496 9673 9505 9707
rect 9505 9673 9539 9707
rect 9539 9673 9548 9707
rect 9496 9664 9548 9673
rect 9588 9664 9640 9716
rect 11152 9664 11204 9716
rect 11520 9664 11572 9716
rect 12348 9664 12400 9716
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6736 9528 6788 9580
rect 7748 9596 7800 9648
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7196 9528 7248 9580
rect 5448 9460 5500 9512
rect 1676 9435 1728 9444
rect 1676 9401 1685 9435
rect 1685 9401 1719 9435
rect 1719 9401 1728 9435
rect 1676 9392 1728 9401
rect 5080 9392 5132 9444
rect 6460 9392 6512 9444
rect 6552 9392 6604 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3148 9324 3200 9376
rect 5908 9324 5960 9376
rect 6276 9324 6328 9376
rect 7196 9392 7248 9444
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7564 9460 7616 9512
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9036 9460 9088 9512
rect 10140 9596 10192 9648
rect 9864 9528 9916 9580
rect 10784 9528 10836 9580
rect 11060 9528 11112 9580
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 9312 9392 9364 9444
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 6920 9324 6972 9376
rect 7656 9324 7708 9376
rect 9772 9324 9824 9376
rect 12532 9392 12584 9444
rect 11980 9324 12032 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 1492 8984 1544 9036
rect 2504 9120 2556 9172
rect 3148 9120 3200 9172
rect 4252 9120 4304 9172
rect 5356 9120 5408 9172
rect 2964 8984 3016 9036
rect 4068 9052 4120 9104
rect 4988 9052 5040 9104
rect 5632 9052 5684 9104
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5264 8916 5316 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6644 9120 6696 9172
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 10324 9163 10376 9172
rect 7196 9120 7248 9129
rect 5356 8916 5408 8925
rect 2320 8891 2372 8900
rect 2320 8857 2329 8891
rect 2329 8857 2363 8891
rect 2363 8857 2372 8891
rect 2320 8848 2372 8857
rect 2504 8780 2556 8832
rect 3056 8780 3108 8832
rect 4712 8848 4764 8900
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6276 8984 6328 9036
rect 7288 8984 7340 9036
rect 7380 8984 7432 9036
rect 9496 9052 9548 9104
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 11152 9120 11204 9172
rect 11888 9120 11940 9172
rect 9864 9052 9916 9061
rect 10232 9052 10284 9104
rect 5724 8848 5776 8900
rect 6736 8916 6788 8968
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 8576 8916 8628 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9220 8926 9272 8978
rect 9588 8993 9597 9006
rect 9597 8993 9631 9006
rect 9631 8993 9640 9006
rect 9588 8954 9640 8993
rect 7196 8891 7248 8900
rect 7196 8857 7205 8891
rect 7205 8857 7239 8891
rect 7239 8857 7248 8891
rect 7196 8848 7248 8857
rect 7564 8848 7616 8900
rect 8944 8891 8996 8900
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 9588 8848 9640 8900
rect 10140 8891 10192 8900
rect 10140 8857 10149 8891
rect 10149 8857 10183 8891
rect 10183 8857 10192 8891
rect 10140 8848 10192 8857
rect 12072 8984 12124 9036
rect 10692 8848 10744 8900
rect 6828 8780 6880 8832
rect 7748 8780 7800 8832
rect 9128 8780 9180 8832
rect 9496 8780 9548 8832
rect 9864 8780 9916 8832
rect 10784 8780 10836 8832
rect 12440 8891 12492 8900
rect 12440 8857 12474 8891
rect 12474 8857 12492 8891
rect 12440 8848 12492 8857
rect 11704 8780 11756 8832
rect 11980 8780 12032 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 2658 8678 2710 8730
rect 2722 8678 2774 8730
rect 2786 8678 2838 8730
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 8658 8678 8710 8730
rect 8722 8678 8774 8730
rect 8786 8678 8838 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 1676 8576 1728 8628
rect 2320 8576 2372 8628
rect 2504 8576 2556 8628
rect 3056 8576 3108 8628
rect 4252 8576 4304 8628
rect 4988 8619 5040 8628
rect 4988 8585 5015 8619
rect 5015 8585 5040 8619
rect 4988 8576 5040 8585
rect 5632 8576 5684 8628
rect 5908 8619 5960 8628
rect 5908 8585 5917 8619
rect 5917 8585 5951 8619
rect 5951 8585 5960 8619
rect 5908 8576 5960 8585
rect 6368 8576 6420 8628
rect 6828 8576 6880 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 2780 8372 2832 8424
rect 2412 8304 2464 8356
rect 5080 8440 5132 8492
rect 5264 8508 5316 8560
rect 5632 8440 5684 8492
rect 7012 8508 7064 8560
rect 10232 8576 10284 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 12440 8576 12492 8628
rect 14004 8508 14056 8560
rect 4068 8372 4120 8424
rect 3516 8304 3568 8356
rect 5816 8372 5868 8424
rect 9128 8440 9180 8492
rect 9496 8440 9548 8492
rect 9772 8440 9824 8492
rect 5724 8304 5776 8356
rect 6828 8304 6880 8356
rect 9312 8372 9364 8424
rect 9588 8372 9640 8424
rect 10324 8440 10376 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 10140 8372 10192 8424
rect 10876 8304 10928 8356
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 4712 8236 4764 8288
rect 7196 8236 7248 8288
rect 8576 8236 8628 8288
rect 9864 8236 9916 8288
rect 11796 8372 11848 8424
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 13544 8440 13596 8492
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 5632 8032 5684 8084
rect 8392 8032 8444 8084
rect 9496 8032 9548 8084
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 2780 7964 2832 8016
rect 3424 7896 3476 7948
rect 4620 7896 4672 7948
rect 1584 7828 1636 7880
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3148 7828 3200 7880
rect 9312 7964 9364 8016
rect 8392 7896 8444 7948
rect 10876 7964 10928 8016
rect 12164 7964 12216 8016
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 9496 7760 9548 7812
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 9128 7692 9180 7744
rect 9220 7692 9272 7744
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 10140 7692 10192 7744
rect 10876 7692 10928 7744
rect 11428 7692 11480 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 8658 7590 8710 7642
rect 8722 7590 8774 7642
rect 8786 7590 8838 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 3148 7488 3200 7540
rect 7012 7488 7064 7540
rect 1676 7352 1728 7404
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 1400 7284 1452 7336
rect 7656 7420 7708 7472
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6920 7352 6972 7404
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 8484 7488 8536 7540
rect 9312 7488 9364 7540
rect 11244 7488 11296 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 9128 7420 9180 7472
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 9220 7352 9272 7404
rect 10048 7420 10100 7472
rect 10140 7352 10192 7404
rect 10692 7352 10744 7404
rect 9496 7284 9548 7336
rect 10876 7216 10928 7268
rect 11980 7352 12032 7404
rect 13452 7352 13504 7404
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 9588 7148 9640 7200
rect 11060 7148 11112 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 11980 7148 12032 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 4068 6944 4120 6996
rect 6828 6944 6880 6996
rect 7104 6944 7156 6996
rect 7656 6944 7708 6996
rect 5908 6876 5960 6928
rect 9220 6876 9272 6928
rect 9588 6944 9640 6996
rect 10048 6944 10100 6996
rect 11704 6876 11756 6928
rect 7564 6808 7616 6860
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5448 6740 5500 6792
rect 6184 6740 6236 6792
rect 6920 6740 6972 6792
rect 7104 6740 7156 6792
rect 9220 6740 9272 6792
rect 8576 6672 8628 6724
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11980 6808 12032 6860
rect 10876 6740 10928 6792
rect 11060 6740 11112 6792
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 7380 6604 7432 6656
rect 9404 6604 9456 6656
rect 9680 6604 9732 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 10692 6604 10744 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11796 6604 11848 6656
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 8658 6502 8710 6554
rect 8722 6502 8774 6554
rect 8786 6502 8838 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 4436 6400 4488 6452
rect 7564 6400 7616 6452
rect 9036 6400 9088 6452
rect 9496 6400 9548 6452
rect 1676 6264 1728 6316
rect 5448 6332 5500 6384
rect 2412 6307 2464 6316
rect 2412 6273 2446 6307
rect 2446 6273 2464 6307
rect 2412 6264 2464 6273
rect 3148 6060 3200 6112
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4068 6264 4120 6316
rect 4160 6264 4212 6316
rect 7840 6332 7892 6384
rect 7196 6264 7248 6316
rect 7748 6264 7800 6316
rect 9312 6332 9364 6384
rect 8668 6264 8720 6316
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 10600 6400 10652 6452
rect 9588 6171 9640 6180
rect 9588 6137 9597 6171
rect 9597 6137 9631 6171
rect 9631 6137 9640 6171
rect 9588 6128 9640 6137
rect 10692 6264 10744 6316
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 10508 6196 10560 6248
rect 8392 6060 8444 6112
rect 8484 6060 8536 6112
rect 9772 6060 9824 6112
rect 9864 6060 9916 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10600 6103 10652 6112
rect 10600 6069 10609 6103
rect 10609 6069 10643 6103
rect 10643 6069 10652 6103
rect 10600 6060 10652 6069
rect 11336 6307 11388 6316
rect 11336 6273 11345 6307
rect 11345 6273 11379 6307
rect 11379 6273 11388 6307
rect 11336 6264 11388 6273
rect 12440 6264 12492 6316
rect 13544 6264 13596 6316
rect 11428 6196 11480 6248
rect 11060 6060 11112 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 2412 5856 2464 5908
rect 4252 5856 4304 5908
rect 5080 5856 5132 5908
rect 5264 5856 5316 5908
rect 5448 5856 5500 5908
rect 4436 5652 4488 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4988 5652 5040 5704
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 8392 5856 8444 5908
rect 9128 5856 9180 5908
rect 11704 5856 11756 5908
rect 13544 5856 13596 5908
rect 10048 5788 10100 5840
rect 10508 5788 10560 5840
rect 12440 5831 12492 5840
rect 12440 5797 12449 5831
rect 12449 5797 12483 5831
rect 12483 5797 12492 5831
rect 12440 5788 12492 5797
rect 7748 5652 7800 5704
rect 8668 5652 8720 5704
rect 9036 5652 9088 5704
rect 9588 5720 9640 5772
rect 4252 5516 4304 5568
rect 4436 5516 4488 5568
rect 5264 5516 5316 5568
rect 8392 5516 8444 5568
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 9864 5652 9916 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 11888 5652 11940 5704
rect 12164 5652 12216 5704
rect 9772 5584 9824 5636
rect 10048 5584 10100 5636
rect 9312 5516 9364 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 8658 5414 8710 5466
rect 8722 5414 8774 5466
rect 8786 5414 8838 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 2412 5244 2464 5296
rect 4252 5312 4304 5364
rect 4620 5312 4672 5364
rect 1676 5176 1728 5228
rect 6000 5244 6052 5296
rect 2320 4972 2372 5024
rect 4068 5176 4120 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 4528 5108 4580 5160
rect 6736 5040 6788 5092
rect 10048 5176 10100 5228
rect 9864 5108 9916 5160
rect 10508 5244 10560 5296
rect 11060 5312 11112 5364
rect 11060 5176 11112 5228
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 5448 4972 5500 5024
rect 7196 4972 7248 5024
rect 10232 4972 10284 5024
rect 10968 5083 11020 5092
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 13084 5244 13136 5296
rect 12072 5176 12124 5228
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 11980 4972 12032 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 4252 4768 4304 4820
rect 7840 4768 7892 4820
rect 8484 4768 8536 4820
rect 9588 4768 9640 4820
rect 8576 4700 8628 4752
rect 3792 4564 3844 4616
rect 4988 4564 5040 4616
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 5448 4607 5500 4616
rect 5448 4573 5482 4607
rect 5482 4573 5500 4607
rect 5448 4564 5500 4573
rect 7380 4564 7432 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 9680 4632 9732 4684
rect 9864 4700 9916 4752
rect 4620 4496 4672 4548
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 7104 4496 7156 4548
rect 7932 4496 7984 4548
rect 8668 4496 8720 4548
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 10600 4632 10652 4684
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 11060 4564 11112 4616
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 11980 4607 12032 4616
rect 11980 4573 12014 4607
rect 12014 4573 12032 4607
rect 11980 4564 12032 4573
rect 11520 4496 11572 4548
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 8658 4326 8710 4378
rect 8722 4326 8774 4378
rect 8786 4326 8838 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 4620 4224 4672 4276
rect 5080 4224 5132 4276
rect 5724 4224 5776 4276
rect 8116 4224 8168 4276
rect 8392 4224 8444 4276
rect 8484 4224 8536 4276
rect 10416 4224 10468 4276
rect 1676 4088 1728 4140
rect 2412 4131 2464 4140
rect 2412 4097 2446 4131
rect 2446 4097 2464 4131
rect 2412 4088 2464 4097
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4988 4088 5040 4140
rect 4528 3952 4580 4004
rect 5356 4020 5408 4072
rect 7840 4156 7892 4208
rect 7932 3952 7984 4004
rect 8392 3952 8444 4004
rect 12164 3952 12216 4004
rect 3608 3884 3660 3936
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 2412 3680 2464 3732
rect 4344 3680 4396 3732
rect 11520 3680 11572 3732
rect 13452 3680 13504 3732
rect 9128 3655 9180 3664
rect 9128 3621 9137 3655
rect 9137 3621 9171 3655
rect 9171 3621 9180 3655
rect 9128 3612 9180 3621
rect 3240 3544 3292 3596
rect 4068 3519 4120 3528
rect 4068 3485 4087 3519
rect 4087 3485 4120 3519
rect 4068 3476 4120 3485
rect 3700 3408 3752 3460
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5172 3544 5224 3596
rect 7380 3544 7432 3596
rect 6000 3476 6052 3528
rect 6920 3476 6972 3528
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 4620 3408 4672 3460
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 6644 3408 6696 3460
rect 6736 3408 6788 3460
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 8576 3408 8628 3460
rect 9036 3476 9088 3528
rect 7012 3340 7064 3392
rect 9588 3340 9640 3392
rect 10784 3408 10836 3460
rect 13360 3408 13412 3460
rect 11060 3340 11112 3392
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 8658 3238 8710 3290
rect 8722 3238 8774 3290
rect 8786 3238 8838 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 4988 3136 5040 3188
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 7748 3136 7800 3188
rect 8300 3136 8352 3188
rect 9128 3136 9180 3188
rect 1676 3000 1728 3052
rect 3056 3043 3108 3052
rect 3056 3009 3090 3043
rect 3090 3009 3108 3043
rect 3056 3000 3108 3009
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 5172 3000 5224 3052
rect 6736 3111 6788 3120
rect 6736 3077 6745 3111
rect 6745 3077 6779 3111
rect 6779 3077 6788 3111
rect 6736 3068 6788 3077
rect 6828 3111 6880 3120
rect 6828 3077 6837 3111
rect 6837 3077 6871 3111
rect 6871 3077 6880 3111
rect 6828 3068 6880 3077
rect 7196 3068 7248 3120
rect 7012 3000 7064 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7932 3000 7984 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 9312 2932 9364 2984
rect 4436 2796 4488 2848
rect 9404 2796 9456 2848
rect 9588 2796 9640 2848
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 3056 2592 3108 2644
rect 4344 2592 4396 2644
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 7104 2592 7156 2644
rect 5264 2524 5316 2576
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 3148 2456 3200 2508
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 4528 2456 4580 2508
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 3884 2388 3936 2440
rect 4436 2388 4488 2440
rect 4804 2388 4856 2440
rect 6000 2388 6052 2440
rect 6920 2456 6972 2508
rect 7012 2456 7064 2508
rect 8576 2388 8628 2440
rect 9404 2388 9456 2440
rect 9496 2388 9548 2440
rect 9864 2388 9916 2440
rect 848 2252 900 2304
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6828 2252 6880 2304
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 11520 2388 11572 2440
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 14004 2388 14056 2440
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 8658 2150 8710 2202
rect 8722 2150 8774 2202
rect 8786 2150 8838 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
<< metal2 >>
rect 846 16364 902 17164
rect 1858 16364 1914 17164
rect 2870 16364 2926 17164
rect 3882 16364 3938 17164
rect 4894 16364 4950 17164
rect 5906 16364 5962 17164
rect 6918 16364 6974 17164
rect 7930 16364 7986 17164
rect 8942 16364 8998 17164
rect 9954 16364 10010 17164
rect 10966 16364 11022 17164
rect 11978 16364 12034 17164
rect 12990 16364 13046 17164
rect 14002 16364 14058 17164
rect 860 14618 888 16364
rect 1872 14906 1900 16364
rect 1780 14878 1900 14906
rect 1780 14618 1808 14878
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2884 14618 2912 16364
rect 3896 14618 3924 16364
rect 4908 14618 4936 16364
rect 5920 14618 5948 16364
rect 6932 14618 6960 16364
rect 7944 14906 7972 16364
rect 7852 14878 7972 14906
rect 7852 14618 7880 14878
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 8956 14618 8984 16364
rect 848 14612 900 14618
rect 848 14554 900 14560
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 10810 1440 13874
rect 1492 13320 1544 13326
rect 1596 13274 1624 13942
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13326 1716 13670
rect 1544 13268 1624 13274
rect 1492 13262 1624 13268
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1504 13246 1624 13262
rect 1596 12850 1624 13246
rect 1780 13002 1808 14350
rect 2656 14172 3032 14181
rect 2712 14170 2736 14172
rect 2792 14170 2816 14172
rect 2872 14170 2896 14172
rect 2952 14170 2976 14172
rect 2712 14118 2722 14170
rect 2966 14118 2976 14170
rect 2712 14116 2736 14118
rect 2792 14116 2816 14118
rect 2872 14116 2896 14118
rect 2952 14116 2976 14118
rect 2656 14107 3032 14116
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 1688 12974 1808 13002
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1688 11778 1716 12974
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1780 12442 1808 12786
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 2424 12442 2452 13874
rect 2656 13084 3032 13093
rect 2712 13082 2736 13084
rect 2792 13082 2816 13084
rect 2872 13082 2896 13084
rect 2952 13082 2976 13084
rect 2712 13030 2722 13082
rect 2966 13030 2976 13082
rect 2712 13028 2736 13030
rect 2792 13028 2816 13030
rect 2872 13028 2896 13030
rect 2952 13028 2976 13030
rect 2656 13019 3032 13028
rect 3068 12986 3096 14350
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3252 14074 3280 14282
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 3068 12374 3096 12922
rect 3344 12918 3372 13126
rect 3436 12986 3464 13874
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 1504 11750 1716 11778
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1504 10690 1532 11750
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 11132 1624 11630
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11354 1716 11494
rect 1780 11354 1808 12174
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1768 11144 1820 11150
rect 1596 11104 1768 11132
rect 1768 11086 1820 11092
rect 1412 10662 1532 10690
rect 1412 7342 1440 10662
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10266 1532 10542
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1780 10130 1808 11086
rect 2332 10674 2360 11630
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11354 2452 11494
rect 2516 11354 2544 12174
rect 2656 11996 3032 12005
rect 2712 11994 2736 11996
rect 2792 11994 2816 11996
rect 2872 11994 2896 11996
rect 2952 11994 2976 11996
rect 2712 11942 2722 11994
rect 2966 11942 2976 11994
rect 2712 11940 2736 11942
rect 2792 11940 2816 11942
rect 2872 11940 2896 11942
rect 2952 11940 2976 11942
rect 2656 11931 3032 11940
rect 3068 11898 3096 12174
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2700 11286 2728 11766
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2688 11280 2740 11286
rect 2792 11257 2820 11698
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2688 11222 2740 11228
rect 2778 11248 2834 11257
rect 2778 11183 2834 11192
rect 2976 11014 3004 11630
rect 3068 11354 3096 11698
rect 3160 11626 3188 12650
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3252 11830 3280 12310
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2656 10908 3032 10917
rect 2712 10906 2736 10908
rect 2792 10906 2816 10908
rect 2872 10906 2896 10908
rect 2952 10906 2976 10908
rect 2712 10854 2722 10906
rect 2966 10854 2976 10906
rect 2712 10852 2736 10854
rect 2792 10852 2816 10854
rect 2872 10852 2896 10854
rect 2952 10852 2976 10854
rect 2656 10843 3032 10852
rect 3160 10810 3188 11562
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2332 10554 2360 10610
rect 2332 10526 2452 10554
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 2332 10266 2360 10406
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1504 9042 1532 10066
rect 2424 9994 2452 10526
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1596 7886 1624 9318
rect 1688 8634 1716 9386
rect 1780 9178 1808 9454
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2424 8974 2452 9930
rect 2516 9178 2544 9998
rect 2792 9926 2820 10610
rect 3068 10266 3096 10678
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2656 9820 3032 9829
rect 2712 9818 2736 9820
rect 2792 9818 2816 9820
rect 2872 9818 2896 9820
rect 2952 9818 2976 9820
rect 2712 9766 2722 9818
rect 2966 9766 2976 9818
rect 2712 9764 2736 9766
rect 2792 9764 2816 9766
rect 2872 9764 2896 9766
rect 2952 9764 2976 9766
rect 2656 9755 3032 9764
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 3068 9058 3096 10202
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2976 9042 3096 9058
rect 2964 9036 3096 9042
rect 3016 9030 3096 9036
rect 2964 8978 3016 8984
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2332 8634 2360 8842
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2424 8362 2452 8910
rect 3068 8838 3096 9030
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2516 8634 2544 8774
rect 2656 8732 3032 8741
rect 2712 8730 2736 8732
rect 2792 8730 2816 8732
rect 2872 8730 2896 8732
rect 2952 8730 2976 8732
rect 2712 8678 2722 8730
rect 2966 8678 2976 8730
rect 2712 8676 2736 8678
rect 2792 8676 2816 8678
rect 2872 8676 2896 8678
rect 2952 8676 2976 8678
rect 2656 8667 3032 8676
rect 3068 8634 3096 8774
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 2792 8022 2820 8366
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 3160 7886 3188 8230
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 1688 7410 1716 7822
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 3160 7546 3188 7686
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1688 6322 1716 7346
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 1688 5234 1716 6258
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 2424 5914 2452 6258
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 4146 1716 5170
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3058 1716 4082
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 2332 2446 2360 4966
rect 2424 4826 2452 5238
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2424 3738 2452 4082
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3068 2650 3096 2994
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2514 3188 6054
rect 3252 3602 3280 11290
rect 3344 11286 3372 12854
rect 3528 12434 3556 14350
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3620 12986 3648 13262
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3436 12406 3556 12434
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3436 7954 3464 12406
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 11558 3556 11834
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11286 3556 11494
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3620 11082 3648 12922
rect 3712 11354 3740 14282
rect 4172 13841 4200 14350
rect 4724 14074 4752 14418
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4158 13832 4214 13841
rect 4158 13767 4214 13776
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3620 9994 3648 10474
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3528 8362 3556 8910
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3620 2446 3648 3878
rect 3712 3466 3740 10542
rect 3804 4622 3832 11698
rect 3896 6322 3924 12854
rect 3988 10606 4016 13466
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12986 4568 13262
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4632 12850 4660 13670
rect 4724 12850 4752 14010
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4908 13462 4936 13874
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 5552 13394 5580 13942
rect 5644 13530 5672 14350
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13734 6224 14214
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 7300 13530 7328 14350
rect 8656 14172 9032 14181
rect 8712 14170 8736 14172
rect 8792 14170 8816 14172
rect 8872 14170 8896 14172
rect 8952 14170 8976 14172
rect 8712 14118 8722 14170
rect 8966 14118 8976 14170
rect 8712 14116 8736 14118
rect 8792 14116 8816 14118
rect 8872 14116 8896 14118
rect 8952 14116 8976 14118
rect 8656 14107 9032 14116
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 7484 13530 7512 13874
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12918 4844 13126
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4632 12753 4660 12786
rect 5000 12782 5028 13262
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12986 5396 13194
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4988 12776 5040 12782
rect 4618 12744 4674 12753
rect 4988 12718 5040 12724
rect 4618 12679 4674 12688
rect 5000 12442 5028 12718
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 11150 4200 11494
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10742 4108 11018
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 4080 9110 4108 10678
rect 4172 10266 4200 11086
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4264 9178 4292 10134
rect 4540 9926 4568 12106
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4632 10470 4660 10950
rect 4724 10470 4752 12310
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4816 11898 4844 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4908 11762 4936 12038
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11150 4844 11494
rect 5092 11354 5120 12786
rect 5460 12782 5488 13262
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4632 10198 4660 10406
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4724 9926 4752 10406
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4540 9722 4568 9862
rect 4632 9722 4660 9862
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4264 8634 4292 9114
rect 4724 8906 4752 9862
rect 4908 9518 4936 9862
rect 5000 9654 5028 11018
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5092 9450 5120 9930
rect 5184 9722 5212 11834
rect 5368 11762 5396 12310
rect 5460 12102 5488 12718
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5552 10470 5580 13330
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5920 12986 5948 13126
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5736 11898 5764 12718
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5828 11898 5856 12650
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5644 11354 5672 11766
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5920 11234 5948 12922
rect 7300 12918 7328 13466
rect 7852 13394 7880 13670
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12986 7420 13262
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 7288 12912 7340 12918
rect 7288 12854 7340 12860
rect 6196 12434 6224 12854
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 5828 11206 5948 11234
rect 5828 11150 5856 11206
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5276 9722 5304 10134
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5368 9586 5396 9862
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5460 9518 5488 9930
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4896 8968 4948 8974
rect 4894 8936 4896 8945
rect 4948 8936 4950 8945
rect 4712 8900 4764 8906
rect 4894 8871 4950 8880
rect 4712 8842 4764 8848
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 4080 8430 4108 8463
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 7206 4108 8366
rect 4724 8294 4752 8842
rect 5000 8634 5028 9046
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5092 8498 5120 9386
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5368 8974 5396 9114
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5276 8566 5304 8910
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4080 7002 4108 7142
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4080 5234 4108 6258
rect 4172 5556 4200 6258
rect 4264 5914 4292 6598
rect 4448 6458 4476 6734
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5574 4476 5646
rect 4252 5568 4304 5574
rect 4172 5528 4252 5556
rect 4252 5510 4304 5516
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4264 5370 4292 5510
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4080 4146 4108 5170
rect 4540 5166 4568 6734
rect 4632 5710 4660 7890
rect 5552 7410 5580 10406
rect 5736 10266 5764 11086
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5736 9874 5764 10202
rect 5828 10062 5856 10202
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5736 9846 5856 9874
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5644 8634 5672 9046
rect 5828 8974 5856 9846
rect 5920 9382 5948 11206
rect 6012 12406 6224 12434
rect 6932 12434 6960 12786
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 6932 12406 7144 12434
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8090 5672 8434
rect 5736 8362 5764 8842
rect 5828 8430 5856 8910
rect 5920 8634 5948 9318
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6934 5948 7346
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5092 5914 5120 6734
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 5914 5304 6598
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4826 4292 4966
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3988 4049 4016 4082
rect 3974 4040 4030 4049
rect 3974 3975 4030 3984
rect 4080 3534 4108 4082
rect 4540 4010 4568 5102
rect 4632 4554 4660 5306
rect 5000 4622 5028 5646
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4632 4282 4660 4490
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3738 4384 3878
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 2446 3924 3334
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4356 2650 4384 2994
rect 4448 2854 4476 3470
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4448 2446 4476 2790
rect 4540 2514 4568 3946
rect 4632 3466 4660 4218
rect 5000 4146 5028 4558
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5092 4282 5120 4422
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3534 5028 4082
rect 5184 3602 5212 4558
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4816 2446 4844 3334
rect 5000 3194 5028 3470
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5184 3058 5212 3538
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5276 2582 5304 5510
rect 5368 4078 5396 6734
rect 5460 6390 5488 6734
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5460 5914 5488 6326
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 6012 5302 6040 12406
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 11830 6316 12106
rect 7116 12102 7144 12406
rect 8404 12238 8432 13670
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12306 8524 13126
rect 8656 13084 9032 13093
rect 8712 13082 8736 13084
rect 8792 13082 8816 13084
rect 8872 13082 8896 13084
rect 8952 13082 8976 13084
rect 8712 13030 8722 13082
rect 8966 13030 8976 13082
rect 8712 13028 8736 13030
rect 8792 13028 8816 13030
rect 8872 13028 8896 13030
rect 8952 13028 8976 13030
rect 8656 13019 9032 13028
rect 9416 13002 9444 13670
rect 9232 12974 9444 13002
rect 9232 12850 9260 12974
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 9220 12844 9272 12850
rect 9404 12844 9456 12850
rect 9220 12786 9272 12792
rect 9324 12804 9404 12832
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8300 12232 8352 12238
rect 8298 12200 8300 12209
rect 8392 12232 8444 12238
rect 8352 12200 8354 12209
rect 8392 12174 8444 12180
rect 8298 12135 8354 12144
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11150 6224 11494
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10266 6224 11086
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 9897 6132 9998
rect 6090 9888 6146 9897
rect 6090 9823 6146 9832
rect 6288 9602 6316 11766
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6368 11348 6420 11354
rect 6420 11308 6500 11336
rect 6368 11290 6420 11296
rect 6472 10266 6500 11308
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6380 10130 6408 10202
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6196 9574 6316 9602
rect 6196 6798 6224 9574
rect 6564 9450 6592 11630
rect 6748 11354 6776 11630
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6656 10062 6684 11018
rect 6748 10674 6776 11086
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6932 10470 6960 11086
rect 7024 10810 7052 11630
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6644 10056 6696 10062
rect 6932 10010 6960 10406
rect 6644 9998 6696 10004
rect 6656 9466 6684 9998
rect 6748 9982 6960 10010
rect 6748 9586 6776 9982
rect 7010 9888 7066 9897
rect 7010 9823 7066 9832
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6552 9444 6604 9450
rect 6656 9438 6776 9466
rect 6552 9386 6604 9392
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 9042 6316 9318
rect 6368 9172 6420 9178
rect 6472 9160 6500 9386
rect 6644 9172 6696 9178
rect 6472 9132 6644 9160
rect 6368 9114 6420 9120
rect 6644 9114 6696 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6380 8634 6408 9114
rect 6748 8974 6776 9438
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6748 8514 6776 8910
rect 6840 8838 6868 9318
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8634 6868 8774
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6748 8486 6868 8514
rect 6840 8362 6868 8486
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6932 7410 6960 9318
rect 7024 8566 7052 9823
rect 7116 9586 7144 12038
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 9586 7236 11086
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9178 7236 9386
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 9042 7328 10202
rect 7392 9994 7420 11290
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7576 10606 7604 11086
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7484 9738 7512 10066
rect 7576 9926 7604 10542
rect 7668 10266 7696 12038
rect 7852 11354 7880 12038
rect 8312 11694 8340 12135
rect 8404 11762 8432 12174
rect 8496 12170 8524 12242
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11898 8524 12106
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8116 11280 8168 11286
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 8114 11248 8116 11257
rect 8168 11248 8170 11257
rect 8114 11183 8170 11192
rect 7760 10674 7788 11183
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7944 10810 7972 10950
rect 8128 10810 8156 10950
rect 8496 10810 8524 11086
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7484 9710 7604 9738
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 9042 7420 9522
rect 7576 9518 7604 9710
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7576 8906 7604 9454
rect 7668 9382 7696 9930
rect 7760 9654 7788 10474
rect 7852 9994 7880 10746
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8974 7696 9318
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7024 7546 7052 8502
rect 7208 8294 7236 8842
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4622 5488 4966
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5736 4282 5764 5170
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 3194 6040 3470
rect 6748 3466 6776 5034
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 6012 2446 6040 3130
rect 6656 2650 6684 3402
rect 6748 3126 6776 3402
rect 6840 3126 6868 6938
rect 6932 6798 6960 7346
rect 7116 7002 7144 7346
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7116 6798 7144 6938
rect 7576 6866 7604 7278
rect 7668 7002 7696 7414
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5914 7236 6258
rect 7392 5914 7420 6598
rect 7576 6458 7604 6802
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7760 6322 7788 8774
rect 7852 8634 7880 9930
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7852 6390 7880 8570
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 8404 8090 8432 10542
rect 8496 10130 8524 10746
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8588 9674 8616 12786
rect 8680 12442 8708 12786
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 8656 11996 9032 12005
rect 8712 11994 8736 11996
rect 8792 11994 8816 11996
rect 8872 11994 8896 11996
rect 8952 11994 8976 11996
rect 8712 11942 8722 11994
rect 8966 11942 8976 11994
rect 8712 11940 8736 11942
rect 8792 11940 8816 11942
rect 8872 11940 8896 11942
rect 8952 11940 8976 11942
rect 8656 11931 9032 11940
rect 9140 11830 9168 12242
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9140 11354 9168 11562
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9232 11234 9260 12786
rect 9324 12374 9352 12804
rect 9404 12786 9456 12792
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9508 12322 9536 13874
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9784 12986 9812 13398
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9600 12424 9628 12718
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9600 12396 9720 12424
rect 9324 11762 9352 12310
rect 9404 12300 9456 12306
rect 9508 12294 9628 12322
rect 9404 12242 9456 12248
rect 9416 12209 9444 12242
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9505 12164 9557 12170
rect 9505 12106 9557 12112
rect 9517 12050 9545 12106
rect 9416 12022 9545 12050
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9140 11218 9260 11234
rect 9128 11212 9260 11218
rect 9180 11206 9260 11212
rect 9128 11154 9180 11160
rect 8656 10908 9032 10917
rect 8712 10906 8736 10908
rect 8792 10906 8816 10908
rect 8872 10906 8896 10908
rect 8952 10906 8976 10908
rect 8712 10854 8722 10906
rect 8966 10854 8976 10906
rect 8712 10852 8736 10854
rect 8792 10852 8816 10854
rect 8872 10852 8896 10854
rect 8952 10852 8976 10854
rect 8656 10843 9032 10852
rect 9232 10810 9260 11206
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9416 10690 9444 12022
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9508 11286 9536 11834
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9140 10662 9444 10690
rect 8956 10198 8984 10610
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8656 9820 9032 9829
rect 8712 9818 8736 9820
rect 8792 9818 8816 9820
rect 8872 9818 8896 9820
rect 8952 9818 8976 9820
rect 8712 9766 8722 9818
rect 8966 9766 8976 9818
rect 8712 9764 8736 9766
rect 8792 9764 8816 9766
rect 8872 9764 8896 9766
rect 8952 9764 8976 9766
rect 8656 9755 9032 9764
rect 8588 9646 9076 9674
rect 9048 9518 9076 9646
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9140 8974 9168 10662
rect 9600 10538 9628 12294
rect 9692 12238 9720 12396
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11830 9720 12174
rect 9784 12170 9812 12650
rect 9876 12306 9904 13806
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9784 11676 9812 12106
rect 9692 11648 9812 11676
rect 9692 11082 9720 11648
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9416 10266 9444 10474
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9508 9722 9536 9998
rect 9600 9722 9628 9998
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9450 9352 9522
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9496 9104 9548 9110
rect 9692 9092 9720 11018
rect 9784 9382 9812 11086
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9586 9904 9998
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9548 9064 9720 9092
rect 9496 9046 9548 9052
rect 9588 9006 9640 9012
rect 9220 8978 9272 8984
rect 8576 8968 8628 8974
rect 9128 8968 9180 8974
rect 8576 8910 8628 8916
rect 8942 8936 8998 8945
rect 8588 8294 8616 8910
rect 9220 8920 9272 8926
rect 9416 8954 9588 8966
rect 9416 8948 9640 8954
rect 9416 8938 9628 8948
rect 9128 8910 9180 8916
rect 8942 8871 8944 8880
rect 8996 8871 8998 8880
rect 8944 8842 8996 8848
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8656 8732 9032 8741
rect 8712 8730 8736 8732
rect 8792 8730 8816 8732
rect 8872 8730 8896 8732
rect 8952 8730 8976 8732
rect 8712 8678 8722 8730
rect 8966 8678 8976 8730
rect 8712 8676 8736 8678
rect 8792 8676 8816 8678
rect 8872 8676 8896 8678
rect 8952 8676 8976 8678
rect 8656 8667 9032 8676
rect 9140 8498 9168 8774
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8404 7954 8432 8026
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8496 7290 8524 7482
rect 8588 7426 8616 8230
rect 9232 7834 9260 8920
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 8022 9352 8366
rect 9416 8294 9444 8938
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8498 9536 8774
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9600 8430 9628 8842
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9416 8266 9536 8294
rect 9508 8090 9536 8266
rect 9692 8090 9720 9064
rect 9784 8498 9812 9318
rect 9876 9110 9904 9522
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9876 8294 9904 8774
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9312 8016 9364 8022
rect 9364 7976 9444 8004
rect 9312 7958 9364 7964
rect 9232 7806 9352 7834
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8656 7644 9032 7653
rect 8712 7642 8736 7644
rect 8792 7642 8816 7644
rect 8872 7642 8896 7644
rect 8952 7642 8976 7644
rect 8712 7590 8722 7642
rect 8966 7590 8976 7642
rect 8712 7588 8736 7590
rect 8792 7588 8816 7590
rect 8872 7588 8896 7590
rect 8952 7588 8976 7590
rect 8656 7579 9032 7588
rect 9140 7478 9168 7686
rect 9128 7472 9180 7478
rect 8588 7398 8708 7426
rect 9128 7414 9180 7420
rect 9232 7410 9260 7686
rect 9324 7546 9352 7806
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 8680 7342 8708 7398
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8668 7336 8720 7342
rect 8496 7262 8616 7290
rect 8668 7278 8720 7284
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8588 6730 8616 7262
rect 9232 6934 9260 7346
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9232 6798 9260 6870
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7760 5710 7788 6258
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8404 5914 8432 6054
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6932 2514 6960 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3058 7052 3334
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7024 2514 7052 2994
rect 7116 2650 7144 4490
rect 7208 3126 7236 4966
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7392 3602 7420 4558
rect 7852 4214 7880 4762
rect 8404 4706 8432 5510
rect 8496 4826 8524 6054
rect 8588 5284 8616 6666
rect 8656 6556 9032 6565
rect 8712 6554 8736 6556
rect 8792 6554 8816 6556
rect 8872 6554 8896 6556
rect 8952 6554 8976 6556
rect 8712 6502 8722 6554
rect 8966 6502 8976 6554
rect 8712 6500 8736 6502
rect 8792 6500 8816 6502
rect 8872 6500 8896 6502
rect 8952 6500 8976 6502
rect 8656 6491 9032 6500
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5710 8708 6258
rect 9048 5710 9076 6394
rect 9232 6322 9260 6734
rect 9324 6390 9352 7482
rect 9416 6662 9444 7976
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 7342 9536 7754
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9508 6458 9536 7278
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 7002 9628 7142
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9140 5642 9168 5850
rect 9508 5760 9536 6394
rect 9600 6186 9628 6938
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9588 5772 9640 5778
rect 9508 5732 9588 5760
rect 9588 5714 9640 5720
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8656 5468 9032 5477
rect 8712 5466 8736 5468
rect 8792 5466 8816 5468
rect 8872 5466 8896 5468
rect 8952 5466 8976 5468
rect 8712 5414 8722 5466
rect 8966 5414 8976 5466
rect 8712 5412 8736 5414
rect 8792 5412 8816 5414
rect 8872 5412 8896 5414
rect 8952 5412 8976 5414
rect 8656 5403 9032 5412
rect 8588 5256 8708 5284
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8312 4678 8432 4706
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7840 4208 7892 4214
rect 7840 4150 7892 4156
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7392 3058 7420 3538
rect 7852 3534 7880 4150
rect 7944 4010 7972 4490
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4282 8156 4422
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8312 4162 8340 4678
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8404 4282 8432 4558
rect 8496 4282 8524 4762
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8312 4134 8432 4162
rect 8404 4010 8432 4134
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 8404 3534 8432 3946
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7760 3194 7788 3470
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7852 3074 7880 3470
rect 8588 3466 8616 4694
rect 8680 4554 8708 5256
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8656 4380 9032 4389
rect 8712 4378 8736 4380
rect 8792 4378 8816 4380
rect 8872 4378 8896 4380
rect 8952 4378 8976 4380
rect 8712 4326 8722 4378
rect 8966 4326 8976 4378
rect 8712 4324 8736 4326
rect 8792 4324 8816 4326
rect 8872 4324 8896 4326
rect 8952 4324 8976 4326
rect 8656 4315 9032 4324
rect 9324 3754 9352 5510
rect 9600 4826 9628 5714
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9692 4690 9720 6598
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9784 5642 9812 6054
rect 9876 5710 9904 6054
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9876 4758 9904 5102
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9048 3726 9352 3754
rect 9048 3534 9076 3726
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8312 3194 8340 3402
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7852 3058 7972 3074
rect 7380 3052 7432 3058
rect 7852 3052 7984 3058
rect 7852 3046 7932 3052
rect 7380 2994 7432 3000
rect 7932 2994 7984 3000
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 8588 2446 8616 3402
rect 8656 3292 9032 3301
rect 8712 3290 8736 3292
rect 8792 3290 8816 3292
rect 8872 3290 8896 3292
rect 8952 3290 8976 3292
rect 8712 3238 8722 3290
rect 8966 3238 8976 3290
rect 8712 3236 8736 3238
rect 8792 3236 8816 3238
rect 8872 3236 8896 3238
rect 8952 3236 8976 3238
rect 8656 3227 9032 3236
rect 9140 3194 9168 3606
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9048 2650 9076 2994
rect 9324 2990 9352 3726
rect 9416 3058 9444 4558
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9416 2938 9444 2994
rect 9416 2910 9536 2938
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9416 2446 9444 2790
rect 9508 2446 9536 2910
rect 9600 2854 9628 3334
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9968 2774 9996 16364
rect 10980 14414 11008 16364
rect 11992 14414 12020 16364
rect 13004 14414 13032 16364
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 11256 13977 11284 14214
rect 11242 13968 11298 13977
rect 10416 13932 10468 13938
rect 11242 13903 11298 13912
rect 10416 13874 10468 13880
rect 10428 13530 10456 13874
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 12646 10088 13262
rect 10244 13190 10272 13398
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 11060 13320 11112 13326
rect 11164 13274 11192 13670
rect 11612 13456 11664 13462
rect 11664 13416 11744 13444
rect 11612 13398 11664 13404
rect 11112 13268 11192 13274
rect 11060 13262 11192 13268
rect 10232 13184 10284 13190
rect 10152 13144 10232 13172
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12238 10088 12582
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10152 12050 10180 13144
rect 10232 13126 10284 13132
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10244 12186 10272 12650
rect 10336 12646 10364 13262
rect 11072 13246 11192 13262
rect 11164 13190 11192 13246
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10796 12986 10824 13126
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10428 12714 10456 12786
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10244 12158 10456 12186
rect 10612 12170 10640 12786
rect 10704 12714 10732 12922
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10428 12102 10456 12158
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10416 12096 10468 12102
rect 10152 12022 10272 12050
rect 10416 12038 10468 12044
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10152 10674 10180 11834
rect 10244 11762 10272 12022
rect 10232 11756 10284 11762
rect 10284 11716 10364 11744
rect 10232 11698 10284 11704
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10060 10198 10088 10542
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10266 10180 10406
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 10152 9654 10180 10202
rect 10244 10062 10272 11154
rect 10336 10810 10364 11716
rect 10428 11558 10456 12038
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10336 10713 10364 10746
rect 10322 10704 10378 10713
rect 10428 10690 10456 11494
rect 10520 11286 10548 11698
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10520 10810 10548 11086
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10428 10662 10548 10690
rect 10322 10639 10378 10648
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 8906 10180 9590
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8430 10180 8842
rect 10244 8634 10272 9046
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10336 8498 10364 9114
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10060 7478 10088 7686
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 7002 10088 7414
rect 10152 7410 10180 7686
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5846 10088 6054
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10428 5710 10456 9930
rect 10520 6798 10548 10662
rect 10612 10606 10640 12106
rect 10704 11762 10732 12650
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 11762 10824 12378
rect 10888 11898 10916 12718
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11072 12238 11100 12378
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11164 12102 11192 13126
rect 11348 12714 11376 13194
rect 11716 13190 11744 13416
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11624 12918 11652 13126
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11532 12442 11560 12786
rect 11716 12764 11744 13126
rect 11808 12850 11836 13738
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11624 12736 11744 12764
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10606 10732 10950
rect 10888 10826 10916 11834
rect 11164 11830 11192 12038
rect 11348 11898 11376 12174
rect 11624 12102 11652 12736
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10796 10798 10916 10826
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10612 10266 10640 10542
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10796 9586 10824 10798
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8634 10732 8842
rect 10796 8838 10824 9522
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10888 8022 10916 8298
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10704 6662 10732 7346
rect 10888 7274 10916 7686
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10888 6798 10916 7210
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10704 6322 10732 6598
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5846 10548 6190
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 5234 10088 5578
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 4622 10088 5170
rect 10244 5030 10272 5510
rect 10520 5302 10548 5782
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10612 4690 10640 6054
rect 10980 5098 11008 11086
rect 11072 10810 11100 11698
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11164 11082 11192 11562
rect 11256 11150 11284 11562
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11244 10736 11296 10742
rect 11058 10704 11114 10713
rect 11244 10678 11296 10684
rect 11058 10639 11114 10648
rect 11072 9586 11100 10639
rect 11256 9994 11284 10678
rect 11532 10606 11560 11018
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11164 9178 11192 9658
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11242 8256 11298 8265
rect 11242 8191 11298 8200
rect 11256 7886 11284 8191
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7546 11284 7822
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6798 11100 7142
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6118 11100 6598
rect 11348 6322 11376 9998
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11440 7750 11468 9862
rect 11532 9722 11560 10542
rect 11624 10266 11652 12038
rect 11716 11558 11744 12174
rect 11808 11762 11836 12786
rect 11992 12646 12020 13126
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11900 12050 11928 12106
rect 11992 12050 12020 12582
rect 11900 12022 12020 12050
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 12176 11694 12204 12650
rect 12164 11688 12216 11694
rect 11992 11648 12164 11676
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10674 11836 10950
rect 11992 10810 12020 11648
rect 12164 11630 12216 11636
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12176 11354 12204 11494
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11716 10266 11744 10610
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11624 9926 11652 10202
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11624 8820 11652 9522
rect 11704 8832 11756 8838
rect 11624 8792 11704 8820
rect 11704 8774 11756 8780
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11440 6254 11468 7686
rect 11716 7206 11744 8774
rect 11808 8430 11836 10610
rect 11992 9674 12020 10746
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12176 10266 12204 10610
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12176 9674 12204 10202
rect 12268 10062 12296 14214
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12360 11898 12388 12106
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11830 12480 12038
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12440 11688 12492 11694
rect 12360 11648 12440 11676
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12360 9722 12388 11648
rect 12440 11630 12492 11636
rect 12544 10810 12572 12106
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11762 12940 12038
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 13004 11626 13032 14214
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 12820 10266 12848 10406
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13556 10198 13584 10406
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 11900 9646 12020 9674
rect 12084 9646 12204 9674
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 11900 9178 11928 9646
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11900 8498 11928 9114
rect 11992 8922 12020 9318
rect 12084 9042 12112 9646
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11992 8894 12112 8922
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8498 12020 8774
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 6934 11744 7142
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6458 11836 6598
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5370 11100 6054
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11716 5574 11744 5850
rect 11900 5710 11928 8434
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 7410 12020 7822
rect 12084 7750 12112 8894
rect 12360 8498 12388 9658
rect 12544 9450 12572 9930
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12452 8634 12480 8842
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 13556 8498 13584 8774
rect 14016 8566 14044 16364
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6866 12020 7142
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5234 11100 5306
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 11716 4622 11744 5510
rect 12084 5234 12112 7686
rect 12176 7546 12204 7958
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12452 5846 12480 6258
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12176 5166 12204 5646
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4622 12020 4966
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4282 10456 4422
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10796 3466 10824 3878
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 11072 3398 11100 4558
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11532 3738 11560 4490
rect 12176 4010 12204 5102
rect 13096 4826 13124 5238
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3058 11100 3334
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 9876 2746 9996 2774
rect 9876 2446 9904 2746
rect 11532 2446 11560 3674
rect 13096 2446 13124 4762
rect 13464 3738 13492 7346
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13556 6322 13584 7278
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 5914 13584 6258
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13372 2650 13400 3402
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 6828 2304 6880 2310
rect 8116 2304 8168 2310
rect 6828 2246 6880 2252
rect 8036 2264 8116 2292
rect 860 800 888 2246
rect 2148 1170 2176 2246
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 3436 1170 3464 2246
rect 4540 1170 4568 2246
rect 5736 1170 5764 2246
rect 2056 1142 2176 1170
rect 3252 1142 3464 1170
rect 4448 1142 4568 1170
rect 5644 1142 5764 1170
rect 2056 800 2084 1142
rect 3252 800 3280 1142
rect 4448 800 4476 1142
rect 5644 800 5672 1142
rect 6840 800 6868 2246
rect 8036 800 8064 2264
rect 9404 2304 9456 2310
rect 8116 2246 8168 2252
rect 9232 2264 9404 2292
rect 8656 2204 9032 2213
rect 8712 2202 8736 2204
rect 8792 2202 8816 2204
rect 8872 2202 8896 2204
rect 8952 2202 8976 2204
rect 8712 2150 8722 2202
rect 8966 2150 8976 2202
rect 8712 2148 8736 2150
rect 8792 2148 8816 2150
rect 8872 2148 8896 2150
rect 8952 2148 8976 2150
rect 8656 2139 9032 2148
rect 9232 800 9260 2264
rect 10508 2304 10560 2310
rect 9404 2246 9456 2252
rect 10428 2264 10508 2292
rect 10428 800 10456 2264
rect 11704 2304 11756 2310
rect 10508 2246 10560 2252
rect 11624 2264 11704 2292
rect 11624 800 11652 2264
rect 12900 2304 12952 2310
rect 11704 2246 11756 2252
rect 12820 2264 12900 2292
rect 12820 800 12848 2264
rect 12900 2246 12952 2252
rect 14016 800 14044 2382
rect 846 0 902 800
rect 2042 0 2098 800
rect 3238 0 3294 800
rect 4434 0 4490 800
rect 5630 0 5686 800
rect 6826 0 6882 800
rect 8022 0 8078 800
rect 9218 0 9274 800
rect 10414 0 10470 800
rect 11610 0 11666 800
rect 12806 0 12862 800
rect 14002 0 14058 800
<< via2 >>
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 2656 14170 2712 14172
rect 2736 14170 2792 14172
rect 2816 14170 2872 14172
rect 2896 14170 2952 14172
rect 2976 14170 3032 14172
rect 2656 14118 2658 14170
rect 2658 14118 2710 14170
rect 2710 14118 2712 14170
rect 2736 14118 2774 14170
rect 2774 14118 2786 14170
rect 2786 14118 2792 14170
rect 2816 14118 2838 14170
rect 2838 14118 2850 14170
rect 2850 14118 2872 14170
rect 2896 14118 2902 14170
rect 2902 14118 2914 14170
rect 2914 14118 2952 14170
rect 2976 14118 2978 14170
rect 2978 14118 3030 14170
rect 3030 14118 3032 14170
rect 2656 14116 2712 14118
rect 2736 14116 2792 14118
rect 2816 14116 2872 14118
rect 2896 14116 2952 14118
rect 2976 14116 3032 14118
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 2656 13082 2712 13084
rect 2736 13082 2792 13084
rect 2816 13082 2872 13084
rect 2896 13082 2952 13084
rect 2976 13082 3032 13084
rect 2656 13030 2658 13082
rect 2658 13030 2710 13082
rect 2710 13030 2712 13082
rect 2736 13030 2774 13082
rect 2774 13030 2786 13082
rect 2786 13030 2792 13082
rect 2816 13030 2838 13082
rect 2838 13030 2850 13082
rect 2850 13030 2872 13082
rect 2896 13030 2902 13082
rect 2902 13030 2914 13082
rect 2914 13030 2952 13082
rect 2976 13030 2978 13082
rect 2978 13030 3030 13082
rect 3030 13030 3032 13082
rect 2656 13028 2712 13030
rect 2736 13028 2792 13030
rect 2816 13028 2872 13030
rect 2896 13028 2952 13030
rect 2976 13028 3032 13030
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 2656 11994 2712 11996
rect 2736 11994 2792 11996
rect 2816 11994 2872 11996
rect 2896 11994 2952 11996
rect 2976 11994 3032 11996
rect 2656 11942 2658 11994
rect 2658 11942 2710 11994
rect 2710 11942 2712 11994
rect 2736 11942 2774 11994
rect 2774 11942 2786 11994
rect 2786 11942 2792 11994
rect 2816 11942 2838 11994
rect 2838 11942 2850 11994
rect 2850 11942 2872 11994
rect 2896 11942 2902 11994
rect 2902 11942 2914 11994
rect 2914 11942 2952 11994
rect 2976 11942 2978 11994
rect 2978 11942 3030 11994
rect 3030 11942 3032 11994
rect 2656 11940 2712 11942
rect 2736 11940 2792 11942
rect 2816 11940 2872 11942
rect 2896 11940 2952 11942
rect 2976 11940 3032 11942
rect 2778 11192 2834 11248
rect 2656 10906 2712 10908
rect 2736 10906 2792 10908
rect 2816 10906 2872 10908
rect 2896 10906 2952 10908
rect 2976 10906 3032 10908
rect 2656 10854 2658 10906
rect 2658 10854 2710 10906
rect 2710 10854 2712 10906
rect 2736 10854 2774 10906
rect 2774 10854 2786 10906
rect 2786 10854 2792 10906
rect 2816 10854 2838 10906
rect 2838 10854 2850 10906
rect 2850 10854 2872 10906
rect 2896 10854 2902 10906
rect 2902 10854 2914 10906
rect 2914 10854 2952 10906
rect 2976 10854 2978 10906
rect 2978 10854 3030 10906
rect 3030 10854 3032 10906
rect 2656 10852 2712 10854
rect 2736 10852 2792 10854
rect 2816 10852 2872 10854
rect 2896 10852 2952 10854
rect 2976 10852 3032 10854
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 2656 9818 2712 9820
rect 2736 9818 2792 9820
rect 2816 9818 2872 9820
rect 2896 9818 2952 9820
rect 2976 9818 3032 9820
rect 2656 9766 2658 9818
rect 2658 9766 2710 9818
rect 2710 9766 2712 9818
rect 2736 9766 2774 9818
rect 2774 9766 2786 9818
rect 2786 9766 2792 9818
rect 2816 9766 2838 9818
rect 2838 9766 2850 9818
rect 2850 9766 2872 9818
rect 2896 9766 2902 9818
rect 2902 9766 2914 9818
rect 2914 9766 2952 9818
rect 2976 9766 2978 9818
rect 2978 9766 3030 9818
rect 3030 9766 3032 9818
rect 2656 9764 2712 9766
rect 2736 9764 2792 9766
rect 2816 9764 2872 9766
rect 2896 9764 2952 9766
rect 2976 9764 3032 9766
rect 2656 8730 2712 8732
rect 2736 8730 2792 8732
rect 2816 8730 2872 8732
rect 2896 8730 2952 8732
rect 2976 8730 3032 8732
rect 2656 8678 2658 8730
rect 2658 8678 2710 8730
rect 2710 8678 2712 8730
rect 2736 8678 2774 8730
rect 2774 8678 2786 8730
rect 2786 8678 2792 8730
rect 2816 8678 2838 8730
rect 2838 8678 2850 8730
rect 2850 8678 2872 8730
rect 2896 8678 2902 8730
rect 2902 8678 2914 8730
rect 2914 8678 2952 8730
rect 2976 8678 2978 8730
rect 2978 8678 3030 8730
rect 3030 8678 3032 8730
rect 2656 8676 2712 8678
rect 2736 8676 2792 8678
rect 2816 8676 2872 8678
rect 2896 8676 2952 8678
rect 2976 8676 3032 8678
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 4158 13776 4214 13832
rect 8656 14170 8712 14172
rect 8736 14170 8792 14172
rect 8816 14170 8872 14172
rect 8896 14170 8952 14172
rect 8976 14170 9032 14172
rect 8656 14118 8658 14170
rect 8658 14118 8710 14170
rect 8710 14118 8712 14170
rect 8736 14118 8774 14170
rect 8774 14118 8786 14170
rect 8786 14118 8792 14170
rect 8816 14118 8838 14170
rect 8838 14118 8850 14170
rect 8850 14118 8872 14170
rect 8896 14118 8902 14170
rect 8902 14118 8914 14170
rect 8914 14118 8952 14170
rect 8976 14118 8978 14170
rect 8978 14118 9030 14170
rect 9030 14118 9032 14170
rect 8656 14116 8712 14118
rect 8736 14116 8792 14118
rect 8816 14116 8872 14118
rect 8896 14116 8952 14118
rect 8976 14116 9032 14118
rect 4618 12688 4674 12744
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 4894 8916 4896 8936
rect 4896 8916 4948 8936
rect 4948 8916 4950 8936
rect 4894 8880 4950 8916
rect 4066 8472 4122 8528
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 3974 3984 4030 4040
rect 8656 13082 8712 13084
rect 8736 13082 8792 13084
rect 8816 13082 8872 13084
rect 8896 13082 8952 13084
rect 8976 13082 9032 13084
rect 8656 13030 8658 13082
rect 8658 13030 8710 13082
rect 8710 13030 8712 13082
rect 8736 13030 8774 13082
rect 8774 13030 8786 13082
rect 8786 13030 8792 13082
rect 8816 13030 8838 13082
rect 8838 13030 8850 13082
rect 8850 13030 8872 13082
rect 8896 13030 8902 13082
rect 8902 13030 8914 13082
rect 8914 13030 8952 13082
rect 8976 13030 8978 13082
rect 8978 13030 9030 13082
rect 9030 13030 9032 13082
rect 8656 13028 8712 13030
rect 8736 13028 8792 13030
rect 8816 13028 8872 13030
rect 8896 13028 8952 13030
rect 8976 13028 9032 13030
rect 8298 12180 8300 12200
rect 8300 12180 8352 12200
rect 8352 12180 8354 12200
rect 8298 12144 8354 12180
rect 6090 9832 6146 9888
rect 7010 9832 7066 9888
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 7746 11192 7802 11248
rect 8114 11228 8116 11248
rect 8116 11228 8168 11248
rect 8168 11228 8170 11248
rect 8114 11192 8170 11228
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 8656 11994 8712 11996
rect 8736 11994 8792 11996
rect 8816 11994 8872 11996
rect 8896 11994 8952 11996
rect 8976 11994 9032 11996
rect 8656 11942 8658 11994
rect 8658 11942 8710 11994
rect 8710 11942 8712 11994
rect 8736 11942 8774 11994
rect 8774 11942 8786 11994
rect 8786 11942 8792 11994
rect 8816 11942 8838 11994
rect 8838 11942 8850 11994
rect 8850 11942 8872 11994
rect 8896 11942 8902 11994
rect 8902 11942 8914 11994
rect 8914 11942 8952 11994
rect 8976 11942 8978 11994
rect 8978 11942 9030 11994
rect 9030 11942 9032 11994
rect 8656 11940 8712 11942
rect 8736 11940 8792 11942
rect 8816 11940 8872 11942
rect 8896 11940 8952 11942
rect 8976 11940 9032 11942
rect 9402 12144 9458 12200
rect 8656 10906 8712 10908
rect 8736 10906 8792 10908
rect 8816 10906 8872 10908
rect 8896 10906 8952 10908
rect 8976 10906 9032 10908
rect 8656 10854 8658 10906
rect 8658 10854 8710 10906
rect 8710 10854 8712 10906
rect 8736 10854 8774 10906
rect 8774 10854 8786 10906
rect 8786 10854 8792 10906
rect 8816 10854 8838 10906
rect 8838 10854 8850 10906
rect 8850 10854 8872 10906
rect 8896 10854 8902 10906
rect 8902 10854 8914 10906
rect 8914 10854 8952 10906
rect 8976 10854 8978 10906
rect 8978 10854 9030 10906
rect 9030 10854 9032 10906
rect 8656 10852 8712 10854
rect 8736 10852 8792 10854
rect 8816 10852 8872 10854
rect 8896 10852 8952 10854
rect 8976 10852 9032 10854
rect 8656 9818 8712 9820
rect 8736 9818 8792 9820
rect 8816 9818 8872 9820
rect 8896 9818 8952 9820
rect 8976 9818 9032 9820
rect 8656 9766 8658 9818
rect 8658 9766 8710 9818
rect 8710 9766 8712 9818
rect 8736 9766 8774 9818
rect 8774 9766 8786 9818
rect 8786 9766 8792 9818
rect 8816 9766 8838 9818
rect 8838 9766 8850 9818
rect 8850 9766 8872 9818
rect 8896 9766 8902 9818
rect 8902 9766 8914 9818
rect 8914 9766 8952 9818
rect 8976 9766 8978 9818
rect 8978 9766 9030 9818
rect 9030 9766 9032 9818
rect 8656 9764 8712 9766
rect 8736 9764 8792 9766
rect 8816 9764 8872 9766
rect 8896 9764 8952 9766
rect 8976 9764 9032 9766
rect 8942 8900 8998 8936
rect 8942 8880 8944 8900
rect 8944 8880 8996 8900
rect 8996 8880 8998 8900
rect 8656 8730 8712 8732
rect 8736 8730 8792 8732
rect 8816 8730 8872 8732
rect 8896 8730 8952 8732
rect 8976 8730 9032 8732
rect 8656 8678 8658 8730
rect 8658 8678 8710 8730
rect 8710 8678 8712 8730
rect 8736 8678 8774 8730
rect 8774 8678 8786 8730
rect 8786 8678 8792 8730
rect 8816 8678 8838 8730
rect 8838 8678 8850 8730
rect 8850 8678 8872 8730
rect 8896 8678 8902 8730
rect 8902 8678 8914 8730
rect 8914 8678 8952 8730
rect 8976 8678 8978 8730
rect 8978 8678 9030 8730
rect 9030 8678 9032 8730
rect 8656 8676 8712 8678
rect 8736 8676 8792 8678
rect 8816 8676 8872 8678
rect 8896 8676 8952 8678
rect 8976 8676 9032 8678
rect 8656 7642 8712 7644
rect 8736 7642 8792 7644
rect 8816 7642 8872 7644
rect 8896 7642 8952 7644
rect 8976 7642 9032 7644
rect 8656 7590 8658 7642
rect 8658 7590 8710 7642
rect 8710 7590 8712 7642
rect 8736 7590 8774 7642
rect 8774 7590 8786 7642
rect 8786 7590 8792 7642
rect 8816 7590 8838 7642
rect 8838 7590 8850 7642
rect 8850 7590 8872 7642
rect 8896 7590 8902 7642
rect 8902 7590 8914 7642
rect 8914 7590 8952 7642
rect 8976 7590 8978 7642
rect 8978 7590 9030 7642
rect 9030 7590 9032 7642
rect 8656 7588 8712 7590
rect 8736 7588 8792 7590
rect 8816 7588 8872 7590
rect 8896 7588 8952 7590
rect 8976 7588 9032 7590
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 8656 6554 8712 6556
rect 8736 6554 8792 6556
rect 8816 6554 8872 6556
rect 8896 6554 8952 6556
rect 8976 6554 9032 6556
rect 8656 6502 8658 6554
rect 8658 6502 8710 6554
rect 8710 6502 8712 6554
rect 8736 6502 8774 6554
rect 8774 6502 8786 6554
rect 8786 6502 8792 6554
rect 8816 6502 8838 6554
rect 8838 6502 8850 6554
rect 8850 6502 8872 6554
rect 8896 6502 8902 6554
rect 8902 6502 8914 6554
rect 8914 6502 8952 6554
rect 8976 6502 8978 6554
rect 8978 6502 9030 6554
rect 9030 6502 9032 6554
rect 8656 6500 8712 6502
rect 8736 6500 8792 6502
rect 8816 6500 8872 6502
rect 8896 6500 8952 6502
rect 8976 6500 9032 6502
rect 8656 5466 8712 5468
rect 8736 5466 8792 5468
rect 8816 5466 8872 5468
rect 8896 5466 8952 5468
rect 8976 5466 9032 5468
rect 8656 5414 8658 5466
rect 8658 5414 8710 5466
rect 8710 5414 8712 5466
rect 8736 5414 8774 5466
rect 8774 5414 8786 5466
rect 8786 5414 8792 5466
rect 8816 5414 8838 5466
rect 8838 5414 8850 5466
rect 8850 5414 8872 5466
rect 8896 5414 8902 5466
rect 8902 5414 8914 5466
rect 8914 5414 8952 5466
rect 8976 5414 8978 5466
rect 8978 5414 9030 5466
rect 9030 5414 9032 5466
rect 8656 5412 8712 5414
rect 8736 5412 8792 5414
rect 8816 5412 8872 5414
rect 8896 5412 8952 5414
rect 8976 5412 9032 5414
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 8656 4378 8712 4380
rect 8736 4378 8792 4380
rect 8816 4378 8872 4380
rect 8896 4378 8952 4380
rect 8976 4378 9032 4380
rect 8656 4326 8658 4378
rect 8658 4326 8710 4378
rect 8710 4326 8712 4378
rect 8736 4326 8774 4378
rect 8774 4326 8786 4378
rect 8786 4326 8792 4378
rect 8816 4326 8838 4378
rect 8838 4326 8850 4378
rect 8850 4326 8872 4378
rect 8896 4326 8902 4378
rect 8902 4326 8914 4378
rect 8914 4326 8952 4378
rect 8976 4326 8978 4378
rect 8978 4326 9030 4378
rect 9030 4326 9032 4378
rect 8656 4324 8712 4326
rect 8736 4324 8792 4326
rect 8816 4324 8872 4326
rect 8896 4324 8952 4326
rect 8976 4324 9032 4326
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 8656 3290 8712 3292
rect 8736 3290 8792 3292
rect 8816 3290 8872 3292
rect 8896 3290 8952 3292
rect 8976 3290 9032 3292
rect 8656 3238 8658 3290
rect 8658 3238 8710 3290
rect 8710 3238 8712 3290
rect 8736 3238 8774 3290
rect 8774 3238 8786 3290
rect 8786 3238 8792 3290
rect 8816 3238 8838 3290
rect 8838 3238 8850 3290
rect 8850 3238 8872 3290
rect 8896 3238 8902 3290
rect 8902 3238 8914 3290
rect 8914 3238 8952 3290
rect 8976 3238 8978 3290
rect 8978 3238 9030 3290
rect 9030 3238 9032 3290
rect 8656 3236 8712 3238
rect 8736 3236 8792 3238
rect 8816 3236 8872 3238
rect 8896 3236 8952 3238
rect 8976 3236 9032 3238
rect 11242 13912 11298 13968
rect 10322 10648 10378 10704
rect 11058 10648 11114 10704
rect 11242 8200 11298 8256
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 8656 2202 8712 2204
rect 8736 2202 8792 2204
rect 8816 2202 8872 2204
rect 8896 2202 8952 2204
rect 8976 2202 9032 2204
rect 8656 2150 8658 2202
rect 8658 2150 8710 2202
rect 8710 2150 8712 2202
rect 8736 2150 8774 2202
rect 8774 2150 8786 2202
rect 8786 2150 8792 2202
rect 8816 2150 8838 2202
rect 8838 2150 8850 2202
rect 8850 2150 8872 2202
rect 8896 2150 8902 2202
rect 8902 2150 8914 2202
rect 8914 2150 8952 2202
rect 8976 2150 8978 2202
rect 8978 2150 9030 2202
rect 9030 2150 9032 2202
rect 8656 2148 8712 2150
rect 8736 2148 8792 2150
rect 8816 2148 8872 2150
rect 8896 2148 8952 2150
rect 8976 2148 9032 2150
<< metal3 >>
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 2646 14176 3042 14177
rect 2646 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3042 14176
rect 2646 14111 3042 14112
rect 8646 14176 9042 14177
rect 8646 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9042 14176
rect 8646 14111 9042 14112
rect 11237 13972 11303 13973
rect 11237 13968 11284 13972
rect 11348 13970 11354 13972
rect 11237 13912 11242 13968
rect 11237 13908 11284 13912
rect 11348 13910 11394 13970
rect 11348 13908 11354 13910
rect 11237 13907 11303 13908
rect 4153 13836 4219 13837
rect 4102 13834 4108 13836
rect 4062 13774 4108 13834
rect 4172 13832 4219 13836
rect 4214 13776 4219 13832
rect 4102 13772 4108 13774
rect 4172 13772 4219 13776
rect 4153 13771 4219 13772
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 2646 13088 3042 13089
rect 2646 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3042 13088
rect 2646 13023 3042 13024
rect 8646 13088 9042 13089
rect 8646 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9042 13088
rect 8646 13023 9042 13024
rect 4613 12748 4679 12749
rect 4613 12746 4660 12748
rect 4568 12744 4660 12746
rect 4568 12688 4618 12744
rect 4568 12686 4660 12688
rect 4613 12684 4660 12686
rect 4724 12684 4730 12748
rect 4613 12683 4679 12684
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 8293 12202 8359 12205
rect 9397 12202 9463 12205
rect 8293 12200 9463 12202
rect 8293 12144 8298 12200
rect 8354 12144 9402 12200
rect 9458 12144 9463 12200
rect 8293 12142 9463 12144
rect 8293 12139 8359 12142
rect 9397 12139 9463 12142
rect 2646 12000 3042 12001
rect 2646 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3042 12000
rect 2646 11935 3042 11936
rect 8646 12000 9042 12001
rect 8646 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9042 12000
rect 8646 11935 9042 11936
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 2773 11250 2839 11253
rect 7741 11250 7807 11253
rect 8109 11250 8175 11253
rect 2773 11248 8175 11250
rect 2773 11192 2778 11248
rect 2834 11192 7746 11248
rect 7802 11192 8114 11248
rect 8170 11192 8175 11248
rect 2773 11190 8175 11192
rect 2773 11187 2839 11190
rect 7741 11187 7807 11190
rect 8109 11187 8175 11190
rect 2646 10912 3042 10913
rect 2646 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3042 10912
rect 2646 10847 3042 10848
rect 8646 10912 9042 10913
rect 8646 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9042 10912
rect 8646 10847 9042 10848
rect 10317 10706 10383 10709
rect 11053 10706 11119 10709
rect 10317 10704 11119 10706
rect 10317 10648 10322 10704
rect 10378 10648 11058 10704
rect 11114 10648 11119 10704
rect 10317 10646 11119 10648
rect 10317 10643 10383 10646
rect 11053 10643 11119 10646
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 6085 9890 6151 9893
rect 7005 9890 7071 9893
rect 6085 9888 7071 9890
rect 6085 9832 6090 9888
rect 6146 9832 7010 9888
rect 7066 9832 7071 9888
rect 6085 9830 7071 9832
rect 6085 9827 6151 9830
rect 7005 9827 7071 9830
rect 2646 9824 3042 9825
rect 2646 9760 2652 9824
rect 2716 9760 2732 9824
rect 2796 9760 2812 9824
rect 2876 9760 2892 9824
rect 2956 9760 2972 9824
rect 3036 9760 3042 9824
rect 2646 9759 3042 9760
rect 8646 9824 9042 9825
rect 8646 9760 8652 9824
rect 8716 9760 8732 9824
rect 8796 9760 8812 9824
rect 8876 9760 8892 9824
rect 8956 9760 8972 9824
rect 9036 9760 9042 9824
rect 8646 9759 9042 9760
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 4889 8938 4955 8941
rect 8937 8938 9003 8941
rect 4889 8936 9003 8938
rect 4889 8880 4894 8936
rect 4950 8880 8942 8936
rect 8998 8880 9003 8936
rect 4889 8878 9003 8880
rect 4889 8875 4955 8878
rect 8937 8875 9003 8878
rect 2646 8736 3042 8737
rect 2646 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3042 8736
rect 2646 8671 3042 8672
rect 8646 8736 9042 8737
rect 8646 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9042 8736
rect 8646 8671 9042 8672
rect 4061 8532 4127 8533
rect 4061 8528 4108 8532
rect 4172 8530 4178 8532
rect 4061 8472 4066 8528
rect 4061 8468 4108 8472
rect 4172 8470 4218 8530
rect 4172 8468 4178 8470
rect 4061 8467 4127 8468
rect 11237 8260 11303 8261
rect 11237 8258 11284 8260
rect 11192 8256 11284 8258
rect 11192 8200 11242 8256
rect 11192 8198 11284 8200
rect 11237 8196 11284 8198
rect 11348 8196 11354 8260
rect 11237 8195 11303 8196
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 8646 7648 9042 7649
rect 8646 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9042 7648
rect 8646 7583 9042 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 8646 6560 9042 6561
rect 8646 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9042 6560
rect 8646 6495 9042 6496
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 8646 5472 9042 5473
rect 8646 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9042 5472
rect 8646 5407 9042 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 8646 4384 9042 4385
rect 8646 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9042 4384
rect 8646 4319 9042 4320
rect 3969 4042 4035 4045
rect 4654 4042 4660 4044
rect 3969 4040 4660 4042
rect 3969 3984 3974 4040
rect 4030 3984 4660 4040
rect 3969 3982 4660 3984
rect 3969 3979 4035 3982
rect 4654 3980 4660 3982
rect 4724 3980 4730 4044
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 8646 3296 9042 3297
rect 8646 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9042 3296
rect 8646 3231 9042 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 8646 2208 9042 2209
rect 8646 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9042 2208
rect 8646 2143 9042 2144
<< via3 >>
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 2652 14172 2716 14176
rect 2652 14116 2656 14172
rect 2656 14116 2712 14172
rect 2712 14116 2716 14172
rect 2652 14112 2716 14116
rect 2732 14172 2796 14176
rect 2732 14116 2736 14172
rect 2736 14116 2792 14172
rect 2792 14116 2796 14172
rect 2732 14112 2796 14116
rect 2812 14172 2876 14176
rect 2812 14116 2816 14172
rect 2816 14116 2872 14172
rect 2872 14116 2876 14172
rect 2812 14112 2876 14116
rect 2892 14172 2956 14176
rect 2892 14116 2896 14172
rect 2896 14116 2952 14172
rect 2952 14116 2956 14172
rect 2892 14112 2956 14116
rect 2972 14172 3036 14176
rect 2972 14116 2976 14172
rect 2976 14116 3032 14172
rect 3032 14116 3036 14172
rect 2972 14112 3036 14116
rect 8652 14172 8716 14176
rect 8652 14116 8656 14172
rect 8656 14116 8712 14172
rect 8712 14116 8716 14172
rect 8652 14112 8716 14116
rect 8732 14172 8796 14176
rect 8732 14116 8736 14172
rect 8736 14116 8792 14172
rect 8792 14116 8796 14172
rect 8732 14112 8796 14116
rect 8812 14172 8876 14176
rect 8812 14116 8816 14172
rect 8816 14116 8872 14172
rect 8872 14116 8876 14172
rect 8812 14112 8876 14116
rect 8892 14172 8956 14176
rect 8892 14116 8896 14172
rect 8896 14116 8952 14172
rect 8952 14116 8956 14172
rect 8892 14112 8956 14116
rect 8972 14172 9036 14176
rect 8972 14116 8976 14172
rect 8976 14116 9032 14172
rect 9032 14116 9036 14172
rect 8972 14112 9036 14116
rect 11284 13968 11348 13972
rect 11284 13912 11298 13968
rect 11298 13912 11348 13968
rect 11284 13908 11348 13912
rect 4108 13832 4172 13836
rect 4108 13776 4158 13832
rect 4158 13776 4172 13832
rect 4108 13772 4172 13776
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 2652 13084 2716 13088
rect 2652 13028 2656 13084
rect 2656 13028 2712 13084
rect 2712 13028 2716 13084
rect 2652 13024 2716 13028
rect 2732 13084 2796 13088
rect 2732 13028 2736 13084
rect 2736 13028 2792 13084
rect 2792 13028 2796 13084
rect 2732 13024 2796 13028
rect 2812 13084 2876 13088
rect 2812 13028 2816 13084
rect 2816 13028 2872 13084
rect 2872 13028 2876 13084
rect 2812 13024 2876 13028
rect 2892 13084 2956 13088
rect 2892 13028 2896 13084
rect 2896 13028 2952 13084
rect 2952 13028 2956 13084
rect 2892 13024 2956 13028
rect 2972 13084 3036 13088
rect 2972 13028 2976 13084
rect 2976 13028 3032 13084
rect 3032 13028 3036 13084
rect 2972 13024 3036 13028
rect 8652 13084 8716 13088
rect 8652 13028 8656 13084
rect 8656 13028 8712 13084
rect 8712 13028 8716 13084
rect 8652 13024 8716 13028
rect 8732 13084 8796 13088
rect 8732 13028 8736 13084
rect 8736 13028 8792 13084
rect 8792 13028 8796 13084
rect 8732 13024 8796 13028
rect 8812 13084 8876 13088
rect 8812 13028 8816 13084
rect 8816 13028 8872 13084
rect 8872 13028 8876 13084
rect 8812 13024 8876 13028
rect 8892 13084 8956 13088
rect 8892 13028 8896 13084
rect 8896 13028 8952 13084
rect 8952 13028 8956 13084
rect 8892 13024 8956 13028
rect 8972 13084 9036 13088
rect 8972 13028 8976 13084
rect 8976 13028 9032 13084
rect 9032 13028 9036 13084
rect 8972 13024 9036 13028
rect 4660 12744 4724 12748
rect 4660 12688 4674 12744
rect 4674 12688 4724 12744
rect 4660 12684 4724 12688
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 2652 11996 2716 12000
rect 2652 11940 2656 11996
rect 2656 11940 2712 11996
rect 2712 11940 2716 11996
rect 2652 11936 2716 11940
rect 2732 11996 2796 12000
rect 2732 11940 2736 11996
rect 2736 11940 2792 11996
rect 2792 11940 2796 11996
rect 2732 11936 2796 11940
rect 2812 11996 2876 12000
rect 2812 11940 2816 11996
rect 2816 11940 2872 11996
rect 2872 11940 2876 11996
rect 2812 11936 2876 11940
rect 2892 11996 2956 12000
rect 2892 11940 2896 11996
rect 2896 11940 2952 11996
rect 2952 11940 2956 11996
rect 2892 11936 2956 11940
rect 2972 11996 3036 12000
rect 2972 11940 2976 11996
rect 2976 11940 3032 11996
rect 3032 11940 3036 11996
rect 2972 11936 3036 11940
rect 8652 11996 8716 12000
rect 8652 11940 8656 11996
rect 8656 11940 8712 11996
rect 8712 11940 8716 11996
rect 8652 11936 8716 11940
rect 8732 11996 8796 12000
rect 8732 11940 8736 11996
rect 8736 11940 8792 11996
rect 8792 11940 8796 11996
rect 8732 11936 8796 11940
rect 8812 11996 8876 12000
rect 8812 11940 8816 11996
rect 8816 11940 8872 11996
rect 8872 11940 8876 11996
rect 8812 11936 8876 11940
rect 8892 11996 8956 12000
rect 8892 11940 8896 11996
rect 8896 11940 8952 11996
rect 8952 11940 8956 11996
rect 8892 11936 8956 11940
rect 8972 11996 9036 12000
rect 8972 11940 8976 11996
rect 8976 11940 9032 11996
rect 9032 11940 9036 11996
rect 8972 11936 9036 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 2652 10908 2716 10912
rect 2652 10852 2656 10908
rect 2656 10852 2712 10908
rect 2712 10852 2716 10908
rect 2652 10848 2716 10852
rect 2732 10908 2796 10912
rect 2732 10852 2736 10908
rect 2736 10852 2792 10908
rect 2792 10852 2796 10908
rect 2732 10848 2796 10852
rect 2812 10908 2876 10912
rect 2812 10852 2816 10908
rect 2816 10852 2872 10908
rect 2872 10852 2876 10908
rect 2812 10848 2876 10852
rect 2892 10908 2956 10912
rect 2892 10852 2896 10908
rect 2896 10852 2952 10908
rect 2952 10852 2956 10908
rect 2892 10848 2956 10852
rect 2972 10908 3036 10912
rect 2972 10852 2976 10908
rect 2976 10852 3032 10908
rect 3032 10852 3036 10908
rect 2972 10848 3036 10852
rect 8652 10908 8716 10912
rect 8652 10852 8656 10908
rect 8656 10852 8712 10908
rect 8712 10852 8716 10908
rect 8652 10848 8716 10852
rect 8732 10908 8796 10912
rect 8732 10852 8736 10908
rect 8736 10852 8792 10908
rect 8792 10852 8796 10908
rect 8732 10848 8796 10852
rect 8812 10908 8876 10912
rect 8812 10852 8816 10908
rect 8816 10852 8872 10908
rect 8872 10852 8876 10908
rect 8812 10848 8876 10852
rect 8892 10908 8956 10912
rect 8892 10852 8896 10908
rect 8896 10852 8952 10908
rect 8952 10852 8956 10908
rect 8892 10848 8956 10852
rect 8972 10908 9036 10912
rect 8972 10852 8976 10908
rect 8976 10852 9032 10908
rect 9032 10852 9036 10908
rect 8972 10848 9036 10852
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 2652 9820 2716 9824
rect 2652 9764 2656 9820
rect 2656 9764 2712 9820
rect 2712 9764 2716 9820
rect 2652 9760 2716 9764
rect 2732 9820 2796 9824
rect 2732 9764 2736 9820
rect 2736 9764 2792 9820
rect 2792 9764 2796 9820
rect 2732 9760 2796 9764
rect 2812 9820 2876 9824
rect 2812 9764 2816 9820
rect 2816 9764 2872 9820
rect 2872 9764 2876 9820
rect 2812 9760 2876 9764
rect 2892 9820 2956 9824
rect 2892 9764 2896 9820
rect 2896 9764 2952 9820
rect 2952 9764 2956 9820
rect 2892 9760 2956 9764
rect 2972 9820 3036 9824
rect 2972 9764 2976 9820
rect 2976 9764 3032 9820
rect 3032 9764 3036 9820
rect 2972 9760 3036 9764
rect 8652 9820 8716 9824
rect 8652 9764 8656 9820
rect 8656 9764 8712 9820
rect 8712 9764 8716 9820
rect 8652 9760 8716 9764
rect 8732 9820 8796 9824
rect 8732 9764 8736 9820
rect 8736 9764 8792 9820
rect 8792 9764 8796 9820
rect 8732 9760 8796 9764
rect 8812 9820 8876 9824
rect 8812 9764 8816 9820
rect 8816 9764 8872 9820
rect 8872 9764 8876 9820
rect 8812 9760 8876 9764
rect 8892 9820 8956 9824
rect 8892 9764 8896 9820
rect 8896 9764 8952 9820
rect 8952 9764 8956 9820
rect 8892 9760 8956 9764
rect 8972 9820 9036 9824
rect 8972 9764 8976 9820
rect 8976 9764 9032 9820
rect 9032 9764 9036 9820
rect 8972 9760 9036 9764
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 2652 8732 2716 8736
rect 2652 8676 2656 8732
rect 2656 8676 2712 8732
rect 2712 8676 2716 8732
rect 2652 8672 2716 8676
rect 2732 8732 2796 8736
rect 2732 8676 2736 8732
rect 2736 8676 2792 8732
rect 2792 8676 2796 8732
rect 2732 8672 2796 8676
rect 2812 8732 2876 8736
rect 2812 8676 2816 8732
rect 2816 8676 2872 8732
rect 2872 8676 2876 8732
rect 2812 8672 2876 8676
rect 2892 8732 2956 8736
rect 2892 8676 2896 8732
rect 2896 8676 2952 8732
rect 2952 8676 2956 8732
rect 2892 8672 2956 8676
rect 2972 8732 3036 8736
rect 2972 8676 2976 8732
rect 2976 8676 3032 8732
rect 3032 8676 3036 8732
rect 2972 8672 3036 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 8732 8732 8796 8736
rect 8732 8676 8736 8732
rect 8736 8676 8792 8732
rect 8792 8676 8796 8732
rect 8732 8672 8796 8676
rect 8812 8732 8876 8736
rect 8812 8676 8816 8732
rect 8816 8676 8872 8732
rect 8872 8676 8876 8732
rect 8812 8672 8876 8676
rect 8892 8732 8956 8736
rect 8892 8676 8896 8732
rect 8896 8676 8952 8732
rect 8952 8676 8956 8732
rect 8892 8672 8956 8676
rect 8972 8732 9036 8736
rect 8972 8676 8976 8732
rect 8976 8676 9032 8732
rect 9032 8676 9036 8732
rect 8972 8672 9036 8676
rect 4108 8528 4172 8532
rect 4108 8472 4122 8528
rect 4122 8472 4172 8528
rect 4108 8468 4172 8472
rect 11284 8256 11348 8260
rect 11284 8200 11298 8256
rect 11298 8200 11348 8256
rect 11284 8196 11348 8200
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 8732 7644 8796 7648
rect 8732 7588 8736 7644
rect 8736 7588 8792 7644
rect 8792 7588 8796 7644
rect 8732 7584 8796 7588
rect 8812 7644 8876 7648
rect 8812 7588 8816 7644
rect 8816 7588 8872 7644
rect 8872 7588 8876 7644
rect 8812 7584 8876 7588
rect 8892 7644 8956 7648
rect 8892 7588 8896 7644
rect 8896 7588 8952 7644
rect 8952 7588 8956 7644
rect 8892 7584 8956 7588
rect 8972 7644 9036 7648
rect 8972 7588 8976 7644
rect 8976 7588 9032 7644
rect 9032 7588 9036 7644
rect 8972 7584 9036 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 8732 6556 8796 6560
rect 8732 6500 8736 6556
rect 8736 6500 8792 6556
rect 8792 6500 8796 6556
rect 8732 6496 8796 6500
rect 8812 6556 8876 6560
rect 8812 6500 8816 6556
rect 8816 6500 8872 6556
rect 8872 6500 8876 6556
rect 8812 6496 8876 6500
rect 8892 6556 8956 6560
rect 8892 6500 8896 6556
rect 8896 6500 8952 6556
rect 8952 6500 8956 6556
rect 8892 6496 8956 6500
rect 8972 6556 9036 6560
rect 8972 6500 8976 6556
rect 8976 6500 9032 6556
rect 9032 6500 9036 6556
rect 8972 6496 9036 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 8732 5468 8796 5472
rect 8732 5412 8736 5468
rect 8736 5412 8792 5468
rect 8792 5412 8796 5468
rect 8732 5408 8796 5412
rect 8812 5468 8876 5472
rect 8812 5412 8816 5468
rect 8816 5412 8872 5468
rect 8872 5412 8876 5468
rect 8812 5408 8876 5412
rect 8892 5468 8956 5472
rect 8892 5412 8896 5468
rect 8896 5412 8952 5468
rect 8952 5412 8956 5468
rect 8892 5408 8956 5412
rect 8972 5468 9036 5472
rect 8972 5412 8976 5468
rect 8976 5412 9032 5468
rect 9032 5412 9036 5468
rect 8972 5408 9036 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 8732 4380 8796 4384
rect 8732 4324 8736 4380
rect 8736 4324 8792 4380
rect 8792 4324 8796 4380
rect 8732 4320 8796 4324
rect 8812 4380 8876 4384
rect 8812 4324 8816 4380
rect 8816 4324 8872 4380
rect 8872 4324 8876 4380
rect 8812 4320 8876 4324
rect 8892 4380 8956 4384
rect 8892 4324 8896 4380
rect 8896 4324 8952 4380
rect 8952 4324 8956 4380
rect 8892 4320 8956 4324
rect 8972 4380 9036 4384
rect 8972 4324 8976 4380
rect 8976 4324 9032 4380
rect 9032 4324 9036 4380
rect 8972 4320 9036 4324
rect 4660 3980 4724 4044
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 8732 3292 8796 3296
rect 8732 3236 8736 3292
rect 8736 3236 8792 3292
rect 8792 3236 8796 3292
rect 8732 3232 8796 3236
rect 8812 3292 8876 3296
rect 8812 3236 8816 3292
rect 8816 3236 8872 3292
rect 8872 3236 8876 3292
rect 8812 3232 8876 3236
rect 8892 3292 8956 3296
rect 8892 3236 8896 3292
rect 8896 3236 8952 3292
rect 8952 3236 8956 3292
rect 8892 3232 8956 3236
rect 8972 3292 9036 3296
rect 8972 3236 8976 3292
rect 8976 3236 9032 3292
rect 9032 3236 9036 3292
rect 8972 3232 9036 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 8732 2204 8796 2208
rect 8732 2148 8736 2204
rect 8736 2148 8792 2204
rect 8792 2148 8796 2204
rect 8732 2144 8796 2148
rect 8812 2204 8876 2208
rect 8812 2148 8816 2204
rect 8816 2148 8872 2204
rect 8872 2148 8876 2204
rect 8812 2144 8876 2148
rect 8892 2204 8956 2208
rect 8892 2148 8896 2204
rect 8896 2148 8952 2204
rect 8952 2148 8956 2204
rect 8892 2144 8956 2148
rect 8972 2204 9036 2208
rect 8972 2148 8976 2204
rect 8976 2148 9032 2204
rect 9032 2148 9036 2204
rect 8972 2144 9036 2148
<< metal4 >>
rect 1904 14720 2304 14736
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9294 2304 10304
rect 1904 9280 1986 9294
rect 2222 9280 2304 9294
rect 1904 9216 1912 9280
rect 1976 9216 1986 9280
rect 2222 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 9058 1986 9216
rect 2222 9058 2304 9216
rect 1904 8192 2304 9058
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 3294 2304 3776
rect 1904 3058 1986 3294
rect 2222 3058 2304 3294
rect 1904 2752 2304 3058
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 2644 14176 3044 14736
rect 2644 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3044 14176
rect 2644 13088 3044 14112
rect 7904 14720 8304 14736
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 4107 13836 4173 13837
rect 4107 13772 4108 13836
rect 4172 13772 4173 13836
rect 4107 13771 4173 13772
rect 2644 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3044 13088
rect 2644 12000 3044 13024
rect 2644 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3044 12000
rect 2644 10912 3044 11936
rect 2644 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3044 10912
rect 2644 10034 3044 10848
rect 2644 9824 2726 10034
rect 2962 9824 3044 10034
rect 2644 9760 2652 9824
rect 2716 9798 2726 9824
rect 2962 9798 2972 9824
rect 2716 9760 2732 9798
rect 2796 9760 2812 9798
rect 2876 9760 2892 9798
rect 2956 9760 2972 9798
rect 3036 9760 3044 9824
rect 2644 8736 3044 9760
rect 2644 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3044 8736
rect 2644 7648 3044 8672
rect 4110 8533 4170 13771
rect 7904 13632 8304 14656
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 4659 12748 4725 12749
rect 4659 12684 4660 12748
rect 4724 12684 4725 12748
rect 4659 12683 4725 12684
rect 4107 8532 4173 8533
rect 4107 8468 4108 8532
rect 4172 8468 4173 8532
rect 4107 8467 4173 8468
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 4034 3044 4320
rect 4662 4045 4722 12683
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9294 8304 10304
rect 7904 9280 7986 9294
rect 8222 9280 8304 9294
rect 7904 9216 7912 9280
rect 7976 9216 7986 9280
rect 8222 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 9058 7986 9216
rect 8222 9058 8304 9216
rect 7904 8192 8304 9058
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 2644 3798 2726 4034
rect 2962 3798 3044 4034
rect 4659 4044 4725 4045
rect 4659 3980 4660 4044
rect 4724 3980 4725 4044
rect 4659 3979 4725 3980
rect 2644 3296 3044 3798
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 2128 3044 2144
rect 7904 3840 8304 4864
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 3294 8304 3776
rect 7904 3058 7986 3294
rect 8222 3058 8304 3294
rect 7904 2752 8304 3058
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 8644 14176 9044 14736
rect 8644 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9044 14176
rect 8644 13088 9044 14112
rect 11283 13972 11349 13973
rect 11283 13908 11284 13972
rect 11348 13908 11349 13972
rect 11283 13907 11349 13908
rect 8644 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9044 13088
rect 8644 12000 9044 13024
rect 8644 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9044 12000
rect 8644 10912 9044 11936
rect 8644 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9044 10912
rect 8644 10034 9044 10848
rect 8644 9824 8726 10034
rect 8962 9824 9044 10034
rect 8644 9760 8652 9824
rect 8716 9798 8726 9824
rect 8962 9798 8972 9824
rect 8716 9760 8732 9798
rect 8796 9760 8812 9798
rect 8876 9760 8892 9798
rect 8956 9760 8972 9798
rect 9036 9760 9044 9824
rect 8644 8736 9044 9760
rect 8644 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9044 8736
rect 8644 7648 9044 8672
rect 11286 8261 11346 13907
rect 11283 8260 11349 8261
rect 11283 8196 11284 8260
rect 11348 8196 11349 8260
rect 11283 8195 11349 8196
rect 8644 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9044 7648
rect 8644 6560 9044 7584
rect 8644 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9044 6560
rect 8644 5472 9044 6496
rect 8644 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9044 5472
rect 8644 4384 9044 5408
rect 8644 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9044 4384
rect 8644 4034 9044 4320
rect 8644 3798 8726 4034
rect 8962 3798 9044 4034
rect 8644 3296 9044 3798
rect 8644 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9044 3296
rect 8644 2208 9044 3232
rect 8644 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9044 2208
rect 8644 2128 9044 2144
<< via4 >>
rect 1986 9280 2222 9294
rect 1986 9216 1992 9280
rect 1992 9216 2056 9280
rect 2056 9216 2072 9280
rect 2072 9216 2136 9280
rect 2136 9216 2152 9280
rect 2152 9216 2216 9280
rect 2216 9216 2222 9280
rect 1986 9058 2222 9216
rect 1986 3058 2222 3294
rect 2726 9824 2962 10034
rect 2726 9798 2732 9824
rect 2732 9798 2796 9824
rect 2796 9798 2812 9824
rect 2812 9798 2876 9824
rect 2876 9798 2892 9824
rect 2892 9798 2956 9824
rect 2956 9798 2962 9824
rect 7986 9280 8222 9294
rect 7986 9216 7992 9280
rect 7992 9216 8056 9280
rect 8056 9216 8072 9280
rect 8072 9216 8136 9280
rect 8136 9216 8152 9280
rect 8152 9216 8216 9280
rect 8216 9216 8222 9280
rect 7986 9058 8222 9216
rect 2726 3798 2962 4034
rect 7986 3058 8222 3294
rect 8726 9824 8962 10034
rect 8726 9798 8732 9824
rect 8732 9798 8796 9824
rect 8796 9798 8812 9824
rect 8812 9798 8876 9824
rect 8876 9798 8892 9824
rect 8892 9798 8956 9824
rect 8956 9798 8962 9824
rect 8726 3798 8962 4034
<< metal5 >>
rect 1056 10034 13940 10116
rect 1056 9798 2726 10034
rect 2962 9798 8726 10034
rect 8962 9798 13940 10034
rect 1056 9716 13940 9798
rect 1056 9294 13940 9376
rect 1056 9058 1986 9294
rect 2222 9058 7986 9294
rect 8222 9058 13940 9294
rect 1056 8976 13940 9058
rect 1056 4034 13940 4116
rect 1056 3798 2726 4034
rect 2962 3798 8726 4034
rect 8962 3798 13940 4034
rect 1056 3716 13940 3798
rect 1056 3294 13940 3376
rect 1056 3058 1986 3294
rect 2222 3058 7986 3294
rect 8222 3058 13940 3294
rect 1056 2976 13940 3058
use sky130_fd_sc_hd__or4bb_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7728 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp 1704896540
transform 1 0 8004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9476 0 -1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11776 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8280 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _203_
timestamp 1704896540
transform -1 0 8832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_2  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10396 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 1704896540
transform -1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _210_
timestamp 1704896540
transform -1 0 11224 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _213_
timestamp 1704896540
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1704896540
transform -1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10120 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _221_
timestamp 1704896540
transform -1 0 6532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _222_
timestamp 1704896540
transform -1 0 7268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp 1704896540
transform -1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _225_
timestamp 1704896540
transform -1 0 6072 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _226_
timestamp 1704896540
transform -1 0 7176 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _227_
timestamp 1704896540
transform -1 0 5612 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _228_
timestamp 1704896540
transform -1 0 6624 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3312 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6440 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _234_
timestamp 1704896540
transform -1 0 5428 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _237_
timestamp 1704896540
transform 1 0 4416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp 1704896540
transform 1 0 4508 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _239_
timestamp 1704896540
transform -1 0 5980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _240_
timestamp 1704896540
transform 1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _241_
timestamp 1704896540
transform -1 0 6256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _242_
timestamp 1704896540
transform -1 0 5888 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _244_
timestamp 1704896540
transform -1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _245_
timestamp 1704896540
transform -1 0 4048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1748 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _248_
timestamp 1704896540
transform -1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _250_
timestamp 1704896540
transform 1 0 4416 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _251_
timestamp 1704896540
transform 1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _252_
timestamp 1704896540
transform -1 0 4968 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1704896540
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _255_
timestamp 1704896540
transform -1 0 5244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _256_
timestamp 1704896540
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _257_
timestamp 1704896540
transform 1 0 3220 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _258_
timestamp 1704896540
transform 1 0 2668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1704896540
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _260_
timestamp 1704896540
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _261_
timestamp 1704896540
transform 1 0 2392 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _262_
timestamp 1704896540
transform 1 0 1472 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1704896540
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1704896540
transform -1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _265_
timestamp 1704896540
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _267_
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _269_
timestamp 1704896540
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1704896540
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1704896540
transform -1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _272_
timestamp 1704896540
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10120 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1704896540
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _275_
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _277_
timestamp 1704896540
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _278_
timestamp 1704896540
transform 1 0 6808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _280_
timestamp 1704896540
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _281_
timestamp 1704896540
transform 1 0 8832 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _282_
timestamp 1704896540
transform 1 0 9108 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _283_
timestamp 1704896540
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _284_
timestamp 1704896540
transform -1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _285_
timestamp 1704896540
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _286_
timestamp 1704896540
transform -1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1704896540
transform 1 0 10028 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1704896540
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _292_
timestamp 1704896540
transform -1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _293_
timestamp 1704896540
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _294_
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _295_
timestamp 1704896540
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _296_
timestamp 1704896540
transform 1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _297_
timestamp 1704896540
transform -1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _298_
timestamp 1704896540
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _299_
timestamp 1704896540
transform -1 0 8464 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _300_
timestamp 1704896540
transform -1 0 7728 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _301_
timestamp 1704896540
transform -1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1704896540
transform -1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1704896540
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _304_
timestamp 1704896540
transform -1 0 10212 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _305_
timestamp 1704896540
transform -1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _306_
timestamp 1704896540
transform -1 0 7268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _308_
timestamp 1704896540
transform -1 0 4692 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1704896540
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _310_
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _311_
timestamp 1704896540
transform -1 0 4692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1704896540
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1704896540
transform 1 0 3680 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _314_
timestamp 1704896540
transform -1 0 4784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _316_
timestamp 1704896540
transform -1 0 4508 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _317_
timestamp 1704896540
transform -1 0 4232 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1704896540
transform 1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _319_
timestamp 1704896540
transform -1 0 5428 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _320_
timestamp 1704896540
transform -1 0 5428 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _321_
timestamp 1704896540
transform -1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _322_
timestamp 1704896540
transform 1 0 6532 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 1704896540
transform -1 0 8004 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1704896540
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _325_
timestamp 1704896540
transform 1 0 4324 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _326_
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1704896540
transform 1 0 6440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _328_
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _329_
timestamp 1704896540
transform 1 0 5244 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp 1704896540
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1704896540
transform -1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9108 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _334_
timestamp 1704896540
transform 1 0 10580 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11224 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _336_
timestamp 1704896540
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12144 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1704896540
transform -1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _339_
timestamp 1704896540
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _340_
timestamp 1704896540
transform -1 0 11868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_1  _341_
timestamp 1704896540
transform 1 0 11868 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1704896540
transform -1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1704896540
transform 1 0 9108 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _344_
timestamp 1704896540
transform 1 0 9936 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _345_
timestamp 1704896540
transform 1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _346_
timestamp 1704896540
transform 1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 1704896540
transform -1 0 12696 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _349_
timestamp 1704896540
transform -1 0 9016 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1704896540
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _352_
timestamp 1704896540
transform 1 0 10672 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _353_
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _354_
timestamp 1704896540
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _356_
timestamp 1704896540
transform -1 0 10580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1704896540
transform -1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _358_
timestamp 1704896540
transform 1 0 9108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _359_
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _360_
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _361_
timestamp 1704896540
transform 1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12052 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _363_
timestamp 1704896540
transform -1 0 12696 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _364_
timestamp 1704896540
transform 1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8096 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _366_
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _367_
timestamp 1704896540
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _368_
timestamp 1704896540
transform -1 0 7636 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _369_
timestamp 1704896540
transform -1 0 5060 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _371_
timestamp 1704896540
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _372_
timestamp 1704896540
transform 1 0 2668 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _373_
timestamp 1704896540
transform -1 0 3680 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _374_
timestamp 1704896540
transform 1 0 1748 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _375_
timestamp 1704896540
transform 1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _376_
timestamp 1704896540
transform 1 0 1472 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1704896540
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3312 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1704896540
transform 1 0 5888 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1704896540
transform 1 0 4784 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1704896540
transform 1 0 2668 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1704896540
transform 1 0 1472 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1704896540
transform -1 0 5612 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1704896540
transform 1 0 7360 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1704896540
transform -1 0 11132 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1704896540
transform 1 0 10580 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1704896540
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1704896540
transform -1 0 8096 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13248 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1704896540
transform 1 0 6072 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1704896540
transform 1 0 2116 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1704896540
transform 1 0 1932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1704896540
transform 1 0 2116 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1704896540
transform 1 0 2760 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1704896540
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1704896540
transform 1 0 6072 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1704896540
transform -1 0 6440 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1704896540
transform 1 0 5152 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1704896540
transform 1 0 12144 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1704896540
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1704896540
transform -1 0 9844 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _404_
timestamp 1704896540
transform 1 0 9844 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _405_
timestamp 1704896540
transform 1 0 12052 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1704896540
transform 1 0 6900 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1704896540
transform 1 0 12144 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1704896540
transform 1 0 1840 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1704896540
transform -1 0 13616 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1704896540
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 6164 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 6256 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_47
timestamp 1704896540
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1704896540
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_66
timestamp 1704896540
transform 1 0 7176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_74
timestamp 1704896540
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79
timestamp 1704896540
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_93
timestamp 1704896540
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 1704896540
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1704896540
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_118
timestamp 1704896540
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1704896540
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_131
timestamp 1704896540
transform 1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_34
timestamp 1704896540
transform 1 0 4232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_66
timestamp 1704896540
transform 1 0 7176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1704896540
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_133
timestamp 1704896540
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18
timestamp 1704896540
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1704896540
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_37
timestamp 1704896540
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_47
timestamp 1704896540
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_75
timestamp 1704896540
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_91
timestamp 1704896540
transform 1 0 9476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_119
timestamp 1704896540
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_40
timestamp 1704896540
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_44
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_50
timestamp 1704896540
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1704896540
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_80
timestamp 1704896540
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_92
timestamp 1704896540
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_96
timestamp 1704896540
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_102
timestamp 1704896540
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1704896540
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_133
timestamp 1704896540
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_11
timestamp 1704896540
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_17
timestamp 1704896540
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1704896540
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_98
timestamp 1704896540
transform 1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_110
timestamp 1704896540
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_114
timestamp 1704896540
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_131
timestamp 1704896540
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_135
timestamp 1704896540
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_25
timestamp 1704896540
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 1704896540
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1704896540
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_71
timestamp 1704896540
transform 1 0 7636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_83
timestamp 1704896540
transform 1 0 8740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_91
timestamp 1704896540
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_102
timestamp 1704896540
transform 1 0 10488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1704896540
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_121
timestamp 1704896540
transform 1 0 12236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_133
timestamp 1704896540
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 1704896540
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_61
timestamp 1704896540
transform 1 0 6716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_72
timestamp 1704896540
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_80
timestamp 1704896540
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_94
timestamp 1704896540
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_124
timestamp 1704896540
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 1704896540
transform 1 0 4232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_73
timestamp 1704896540
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_84
timestamp 1704896540
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1704896540
transform 1 0 10120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_102
timestamp 1704896540
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_132
timestamp 1704896540
transform 1 0 13248 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1704896540
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_39
timestamp 1704896540
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_70
timestamp 1704896540
transform 1 0 7544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 1704896540
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_93
timestamp 1704896540
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_101
timestamp 1704896540
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_105
timestamp 1704896540
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_110
timestamp 1704896540
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 1704896540
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_134
timestamp 1704896540
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1704896540
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_91
timestamp 1704896540
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1704896540
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1704896540
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_73
timestamp 1704896540
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1704896540
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_91
timestamp 1704896540
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_101
timestamp 1704896540
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_107
timestamp 1704896540
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_133
timestamp 1704896540
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_9
timestamp 1704896540
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1704896540
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_45
timestamp 1704896540
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_65
timestamp 1704896540
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_90
timestamp 1704896540
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_98
timestamp 1704896540
transform 1 0 10120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1704896540
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_124
timestamp 1704896540
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_129
timestamp 1704896540
transform 1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_135
timestamp 1704896540
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_36
timestamp 1704896540
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_59
timestamp 1704896540
transform 1 0 6532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_67
timestamp 1704896540
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_75
timestamp 1704896540
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_117
timestamp 1704896540
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_11
timestamp 1704896540
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_23
timestamp 1704896540
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_35
timestamp 1704896540
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_47
timestamp 1704896540
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_90
timestamp 1704896540
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_94
timestamp 1704896540
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1704896540
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_118
timestamp 1704896540
transform 1 0 11960 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_130
timestamp 1704896540
transform 1 0 13064 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_43
timestamp 1704896540
transform 1 0 5060 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_66
timestamp 1704896540
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1704896540
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_92
timestamp 1704896540
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_132
timestamp 1704896540
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_17
timestamp 1704896540
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_24
timestamp 1704896540
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_61
timestamp 1704896540
transform 1 0 6716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_75
timestamp 1704896540
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_94
timestamp 1704896540
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_102
timestamp 1704896540
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1704896540
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_10
timestamp 1704896540
transform 1 0 2024 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1704896540
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_35
timestamp 1704896540
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_43
timestamp 1704896540
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_47
timestamp 1704896540
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_68
timestamp 1704896540
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_72
timestamp 1704896540
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1704896540
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_90
timestamp 1704896540
transform 1 0 9384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_101
timestamp 1704896540
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_110
timestamp 1704896540
transform 1 0 11224 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_122
timestamp 1704896540
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_134
timestamp 1704896540
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_26
timestamp 1704896540
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_32
timestamp 1704896540
transform 1 0 4048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_36
timestamp 1704896540
transform 1 0 4416 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7084 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_78
timestamp 1704896540
transform 1 0 8280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_86
timestamp 1704896540
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_94
timestamp 1704896540
transform 1 0 9752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_103
timestamp 1704896540
transform 1 0 10580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1704896540
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_129
timestamp 1704896540
transform 1 0 12972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_135
timestamp 1704896540
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1704896540
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_11
timestamp 1704896540
transform 1 0 2116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_20
timestamp 1704896540
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_35
timestamp 1704896540
transform 1 0 4324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_43
timestamp 1704896540
transform 1 0 5060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_55
timestamp 1704896540
transform 1 0 6164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_64
timestamp 1704896540
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 1704896540
transform 1 0 7360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1704896540
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_92
timestamp 1704896540
transform 1 0 9568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_96
timestamp 1704896540
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_31
timestamp 1704896540
transform 1 0 3956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_37
timestamp 1704896540
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_42
timestamp 1704896540
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 1704896540
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_68
timestamp 1704896540
transform 1 0 7360 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_83
timestamp 1704896540
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_91
timestamp 1704896540
transform 1 0 9476 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_97
timestamp 1704896540
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 1704896540
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_121
timestamp 1704896540
transform 1 0 12236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_133
timestamp 1704896540
transform 1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1704896540
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_42
timestamp 1704896540
transform 1 0 4968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_50
timestamp 1704896540
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_71
timestamp 1704896540
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1704896540
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_92
timestamp 1704896540
transform 1 0 9568 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_119
timestamp 1704896540
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_131
timestamp 1704896540
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_135
timestamp 1704896540
transform 1 0 13524 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_133
timestamp 1704896540
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_6
timestamp 1704896540
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_12
timestamp 1704896540
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 1704896540
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_34
timestamp 1704896540
transform 1 0 4232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_45
timestamp 1704896540
transform 1 0 5244 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_57
timestamp 1704896540
transform 1 0 6348 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_63
timestamp 1704896540
transform 1 0 6900 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_67
timestamp 1704896540
transform 1 0 7268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_78
timestamp 1704896540
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_89
timestamp 1704896540
transform 1 0 9292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_101
timestamp 1704896540
transform 1 0 10396 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_107
timestamp 1704896540
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_111
timestamp 1704896540
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_113
timestamp 1704896540
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_122
timestamp 1704896540
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_133
timestamp 1704896540
transform 1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1704896540
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1704896540
transform -1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1704896540
transform -1 0 3680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1704896540
transform -1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1704896540
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1704896540
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output13
timestamp 1704896540
transform -1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 1704896540
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 1704896540
transform -1 0 9292 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output16
timestamp 1704896540
transform -1 0 8280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1704896540
transform 1 0 6992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 1704896540
transform -1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp 1704896540
transform -1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1704896540
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1704896540
transform 1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output22
timestamp 1704896540
transform -1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output24
timestamp 1704896540
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 13892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 13892 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 13892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 13892 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 13892 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 13892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 13892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 13892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 13892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 13892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_64
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_66
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_67
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_68
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_69
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_70
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_71
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_72
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_73
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_74
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_75
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_76
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_77
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_78
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_79
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_81
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_82
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_83
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_84
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_85
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_86
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_87
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_88
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_89
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_92
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_93
timestamp 1704896540
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_94
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_95
timestamp 1704896540
transform 1 0 11408 0 1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 2644 2128 3044 14736 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8644 2128 9044 14736 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3716 13940 4116 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9716 13940 10116 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1904 2128 2304 14736 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7904 2128 8304 14736 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2976 13940 3376 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8976 13940 9376 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 analog_comparator_out
port 2 nsew signal input
flabel metal2 s 11978 16364 12034 17164 0 FreeSans 224 90 0 0 calib_enable
port 3 nsew signal input
flabel metal2 s 14002 16364 14058 17164 0 FreeSans 224 90 0 0 clk
port 4 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 comparator_nen
port 5 nsew signal tristate
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 dac_set[0]
port 6 nsew signal tristate
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 dac_set[1]
port 7 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 dac_set[2]
port 8 nsew signal tristate
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 dac_set[3]
port 9 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 dac_set[4]
port 10 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 dac_set[5]
port 11 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 dac_set[6]
port 12 nsew signal tristate
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 dac_set[7]
port 13 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 do_calibrate
port 14 nsew signal tristate
flabel metal2 s 8942 16364 8998 17164 0 FreeSans 224 90 0 0 result[0]
port 15 nsew signal tristate
flabel metal2 s 7930 16364 7986 17164 0 FreeSans 224 90 0 0 result[1]
port 16 nsew signal tristate
flabel metal2 s 6918 16364 6974 17164 0 FreeSans 224 90 0 0 result[2]
port 17 nsew signal tristate
flabel metal2 s 5906 16364 5962 17164 0 FreeSans 224 90 0 0 result[3]
port 18 nsew signal tristate
flabel metal2 s 4894 16364 4950 17164 0 FreeSans 224 90 0 0 result[4]
port 19 nsew signal tristate
flabel metal2 s 3882 16364 3938 17164 0 FreeSans 224 90 0 0 result[5]
port 20 nsew signal tristate
flabel metal2 s 2870 16364 2926 17164 0 FreeSans 224 90 0 0 result[6]
port 21 nsew signal tristate
flabel metal2 s 1858 16364 1914 17164 0 FreeSans 224 90 0 0 result[7]
port 22 nsew signal tristate
flabel metal2 s 846 16364 902 17164 0 FreeSans 224 90 0 0 result_ready
port 23 nsew signal tristate
flabel metal2 s 12990 16364 13046 17164 0 FreeSans 224 90 0 0 rst
port 24 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 thresh_sel
port 25 nsew signal tristate
flabel metal2 s 9954 16364 10010 17164 0 FreeSans 224 90 0 0 use_ext_thresh
port 26 nsew signal input
flabel metal2 s 10966 16364 11022 17164 0 FreeSans 224 90 0 0 user_enable
port 27 nsew signal input
rlabel metal1 7498 14144 7498 14144 0 VGND
rlabel metal1 7498 14688 7498 14688 0 VPWR
rlabel metal2 3450 13430 3450 13430 0 _000_
rlabel metal2 5382 13090 5382 13090 0 _001_
rlabel metal1 1778 7786 1778 7786 0 _002_
rlabel metal1 4692 13430 4692 13430 0 _003_
rlabel metal1 3077 7446 3077 7446 0 _004_
rlabel metal1 1840 12410 1840 12410 0 _005_
rlabel metal1 5489 7446 5489 7446 0 _006_
rlabel metal1 7999 3094 7999 3094 0 _007_
rlabel metal1 10216 3026 10216 3026 0 _008_
rlabel viali 10897 3502 10897 3502 0 _009_
rlabel via1 12001 4590 12001 4590 0 _010_
rlabel metal1 8050 3978 8050 3978 0 _011_
rlabel metal2 7222 6086 7222 6086 0 _012_
rlabel metal2 12466 6052 12466 6052 0 _013_
rlabel metal1 6532 7378 6532 7378 0 _014_
rlabel metal1 2530 5882 2530 5882 0 _015_
rlabel metal2 2438 5032 2438 5032 0 _016_
rlabel metal1 2484 3706 2484 3706 0 _017_
rlabel metal1 3128 2618 3128 2618 0 _018_
rlabel metal1 4820 3026 4820 3026 0 _019_
rlabel metal1 6527 3434 6527 3434 0 _020_
rlabel metal1 6317 5610 6317 5610 0 _021_
rlabel via1 5469 4590 5469 4590 0 _022_
rlabel metal1 12098 10540 12098 10540 0 _023_
rlabel metal2 12466 8738 12466 8738 0 _024_
rlabel via1 9526 13906 9526 13906 0 _025_
rlabel metal1 10488 13498 10488 13498 0 _026_
rlabel metal1 12190 11832 12190 11832 0 _027_
rlabel metal1 7544 13498 7544 13498 0 _028_
rlabel metal1 2576 12410 2576 12410 0 _029_
rlabel via1 1697 13294 1697 13294 0 _030_
rlabel metal1 5060 9962 5060 9962 0 _031_
rlabel metal1 4140 10166 4140 10166 0 _032_
rlabel metal1 6486 9962 6486 9962 0 _033_
rlabel metal2 5382 9724 5382 9724 0 _034_
rlabel metal1 5244 9554 5244 9554 0 _035_
rlabel metal1 4738 9486 4738 9486 0 _036_
rlabel metal1 4278 9894 4278 9894 0 _037_
rlabel metal1 2254 8874 2254 8874 0 _038_
rlabel metal1 2714 11628 2714 11628 0 _039_
rlabel metal1 3611 12682 3611 12682 0 _040_
rlabel metal1 1886 10098 1886 10098 0 _041_
rlabel metal2 5014 10336 5014 10336 0 _042_
rlabel metal1 7268 9554 7268 9554 0 _043_
rlabel metal1 5106 11118 5106 11118 0 _044_
rlabel metal1 4968 12886 4968 12886 0 _045_
rlabel metal1 5060 9690 5060 9690 0 _046_
rlabel metal1 5612 11798 5612 11798 0 _047_
rlabel metal1 5796 12818 5796 12818 0 _048_
rlabel metal1 5842 12614 5842 12614 0 _049_
rlabel metal1 2346 8534 2346 8534 0 _050_
rlabel metal1 4278 11730 4278 11730 0 _051_
rlabel metal1 2622 11594 2622 11594 0 _052_
rlabel metal2 1794 9316 1794 9316 0 _053_
rlabel metal1 1886 8602 1886 8602 0 _054_
rlabel metal1 1518 7854 1518 7854 0 _055_
rlabel metal1 4968 12818 4968 12818 0 _056_
rlabel metal1 4649 12954 4649 12954 0 _057_
rlabel metal1 6946 8058 6946 8058 0 _058_
rlabel via1 5006 8602 5006 8602 0 _059_
rlabel metal1 3450 8364 3450 8364 0 _060_
rlabel metal1 2622 8534 2622 8534 0 _061_
rlabel metal1 3174 8330 3174 8330 0 _062_
rlabel metal1 3266 7854 3266 7854 0 _063_
rlabel metal1 1610 11186 1610 11186 0 _064_
rlabel metal1 2162 11254 2162 11254 0 _065_
rlabel metal1 1886 11322 1886 11322 0 _066_
rlabel metal2 5382 5406 5382 5406 0 _067_
rlabel metal1 4784 2482 4784 2482 0 _068_
rlabel metal1 11362 7378 11362 7378 0 _069_
rlabel metal1 9246 13226 9246 13226 0 _070_
rlabel metal1 8970 3468 8970 3468 0 _071_
rlabel metal1 10994 5134 10994 5134 0 _072_
rlabel metal1 10020 5270 10020 5270 0 _073_
rlabel metal1 8832 2414 8832 2414 0 _074_
rlabel metal1 9614 5678 9614 5678 0 _075_
rlabel metal1 8234 5712 8234 5712 0 _076_
rlabel metal1 9108 3502 9108 3502 0 _077_
rlabel metal1 8832 3638 8832 3638 0 _078_
rlabel metal1 7406 13328 7406 13328 0 _079_
rlabel metal2 9062 2822 9062 2822 0 _080_
rlabel metal1 10488 11730 10488 11730 0 _081_
rlabel metal1 10350 12682 10350 12682 0 _082_
rlabel metal1 10718 6800 10718 6800 0 _083_
rlabel metal1 10166 6630 10166 6630 0 _084_
rlabel metal1 10961 5338 10961 5338 0 _085_
rlabel metal1 10810 4658 10810 4658 0 _086_
rlabel metal1 10258 4148 10258 4148 0 _087_
rlabel metal1 10534 4114 10534 4114 0 _088_
rlabel metal1 12006 5168 12006 5168 0 _089_
rlabel metal1 11868 5202 11868 5202 0 _090_
rlabel metal1 8418 4624 8418 4624 0 _091_
rlabel metal1 7912 6290 7912 6290 0 _092_
rlabel metal1 8418 4794 8418 4794 0 _093_
rlabel metal1 8142 4182 8142 4182 0 _094_
rlabel metal1 7774 5542 7774 5542 0 _095_
rlabel viali 12472 5678 12472 5678 0 _096_
rlabel metal1 10120 4998 10120 4998 0 _097_
rlabel metal1 8694 5202 8694 5202 0 _098_
rlabel metal1 7314 4998 7314 4998 0 _099_
rlabel metal1 5198 3400 5198 3400 0 _100_
rlabel metal1 4324 6426 4324 6426 0 _101_
rlabel metal1 2806 5746 2806 5746 0 _102_
rlabel metal1 4324 5202 4324 5202 0 _103_
rlabel metal1 2691 4590 2691 4590 0 _104_
rlabel metal1 4416 4114 4416 4114 0 _105_
rlabel metal1 2714 3604 2714 3604 0 _106_
rlabel metal1 3956 2414 3956 2414 0 _107_
rlabel metal1 3358 2448 3358 2448 0 _108_
rlabel metal1 5014 2414 5014 2414 0 _109_
rlabel metal1 4692 2618 4692 2618 0 _110_
rlabel metal1 7452 3162 7452 3162 0 _111_
rlabel metal1 6854 2448 6854 2448 0 _112_
rlabel metal1 5014 5882 5014 5882 0 _113_
rlabel metal1 5980 5678 5980 5678 0 _114_
rlabel metal1 5290 4114 5290 4114 0 _115_
rlabel metal1 5704 4250 5704 4250 0 _116_
rlabel metal1 12926 10064 12926 10064 0 _117_
rlabel metal1 12604 9962 12604 9962 0 _118_
rlabel metal1 12650 11696 12650 11696 0 _119_
rlabel metal2 10994 8092 10994 8092 0 _120_
rlabel metal2 11822 9520 11822 9520 0 _121_
rlabel metal2 12834 10336 12834 10336 0 _122_
rlabel metal1 12282 8432 12282 8432 0 _123_
rlabel metal1 11040 9010 11040 9010 0 _124_
rlabel metal2 12006 8636 12006 8636 0 _125_
rlabel metal1 8556 10710 8556 10710 0 _126_
rlabel metal1 9476 10234 9476 10234 0 _127_
rlabel via1 10628 12818 10628 12818 0 _128_
rlabel metal1 10580 10642 10580 10642 0 _129_
rlabel metal1 9522 10608 9522 10608 0 _130_
rlabel metal1 9430 13260 9430 13260 0 _131_
rlabel metal1 8878 10676 8878 10676 0 _132_
rlabel metal1 11224 12886 11224 12886 0 _133_
rlabel metal2 10810 13056 10810 13056 0 _134_
rlabel metal1 11316 12410 11316 12410 0 _135_
rlabel metal1 11960 12614 11960 12614 0 _136_
rlabel metal1 11270 13362 11270 13362 0 _137_
rlabel metal1 10580 13294 10580 13294 0 _138_
rlabel metal1 12696 11798 12696 11798 0 _139_
rlabel metal1 9752 12614 9752 12614 0 _140_
rlabel metal2 10810 12070 10810 12070 0 _141_
rlabel metal1 11270 11662 11270 11662 0 _142_
rlabel metal1 11178 11866 11178 11866 0 _143_
rlabel metal1 12420 11730 12420 11730 0 _144_
rlabel metal2 8602 11239 8602 11239 0 _145_
rlabel metal1 8096 12954 8096 12954 0 _146_
rlabel metal1 8694 13362 8694 13362 0 _147_
rlabel metal1 7728 13294 7728 13294 0 _148_
rlabel metal1 3818 11118 3818 11118 0 _149_
rlabel metal1 3128 11866 3128 11866 0 _150_
rlabel metal2 2530 11764 2530 11764 0 _151_
rlabel metal1 2392 10098 2392 10098 0 _152_
rlabel metal1 1656 10234 1656 10234 0 _153_
rlabel metal1 1978 10506 1978 10506 0 _154_
rlabel metal1 1702 10778 1702 10778 0 _155_
rlabel metal1 6762 8500 6762 8500 0 _156_
rlabel metal1 2300 10030 2300 10030 0 _157_
rlabel metal1 7866 11220 7866 11220 0 _158_
rlabel metal1 10994 7310 10994 7310 0 _159_
rlabel metal1 10442 5236 10442 5236 0 _160_
rlabel metal1 11316 12750 11316 12750 0 _161_
rlabel metal1 6716 10438 6716 10438 0 _162_
rlabel metal1 11362 7786 11362 7786 0 _163_
rlabel metal1 8326 7922 8326 7922 0 _164_
rlabel metal1 11408 7718 11408 7718 0 _165_
rlabel metal1 6854 10778 6854 10778 0 _166_
rlabel metal1 10810 8976 10810 8976 0 _167_
rlabel metal1 6118 11118 6118 11118 0 _168_
rlabel metal1 6624 11322 6624 11322 0 _169_
rlabel metal1 10074 4794 10074 4794 0 _170_
rlabel metal1 7958 9044 7958 9044 0 _171_
rlabel metal1 2806 11798 2806 11798 0 _172_
rlabel metal1 11914 12818 11914 12818 0 _173_
rlabel metal1 7958 10710 7958 10710 0 _174_
rlabel metal1 7682 10608 7682 10608 0 _175_
rlabel metal1 6026 11730 6026 11730 0 _176_
rlabel metal1 6946 9452 6946 9452 0 _177_
rlabel via1 6565 11662 6565 11662 0 _178_
rlabel metal1 3956 12818 3956 12818 0 _179_
rlabel metal1 7406 10234 7406 10234 0 _180_
rlabel metal1 5336 8534 5336 8534 0 _181_
rlabel metal1 9476 7514 9476 7514 0 _182_
rlabel metal1 9200 8874 9200 8874 0 _183_
rlabel metal2 9292 10676 9292 10676 0 _184_
rlabel via2 4922 8925 4922 8925 0 _185_
rlabel metal1 4278 11050 4278 11050 0 _186_
rlabel metal1 9752 8466 9752 8466 0 _187_
rlabel metal1 5934 8908 5934 8908 0 _188_
rlabel metal2 14030 1588 14030 1588 0 analog_comparator_out
rlabel metal1 12052 14382 12052 14382 0 calib_enable
rlabel metal2 14030 12454 14030 12454 0 clk
rlabel metal2 10442 7820 10442 7820 0 clknet_0_clk
rlabel metal1 1932 6290 1932 6290 0 clknet_2_0__leaf_clk
rlabel metal1 1886 13940 1886 13940 0 clknet_2_1__leaf_clk
rlabel metal1 13386 6290 13386 6290 0 clknet_2_2__leaf_clk
rlabel metal1 12144 9010 12144 9010 0 clknet_2_3__leaf_clk
rlabel metal2 12834 1520 12834 1520 0 comparator_nen
rlabel metal2 874 1520 874 1520 0 dac_set[0]
rlabel metal2 2070 959 2070 959 0 dac_set[1]
rlabel metal2 3266 959 3266 959 0 dac_set[2]
rlabel metal2 4462 959 4462 959 0 dac_set[3]
rlabel metal2 5658 959 5658 959 0 dac_set[4]
rlabel metal2 6854 1520 6854 1520 0 dac_set[5]
rlabel metal2 8050 1520 8050 1520 0 dac_set[6]
rlabel metal2 9246 1520 9246 1520 0 dac_set[7]
rlabel metal2 11638 1520 11638 1520 0 do_calibrate
rlabel metal2 13386 3026 13386 3026 0 net1
rlabel metal1 5980 2414 5980 2414 0 net10
rlabel metal1 7084 2414 7084 2414 0 net11
rlabel metal1 8326 2482 8326 2482 0 net12
rlabel metal1 6578 4488 6578 4488 0 net13
rlabel metal1 11730 2414 11730 2414 0 net14
rlabel metal2 4738 14246 4738 14246 0 net15
rlabel metal2 7314 13940 7314 13940 0 net16
rlabel metal2 4646 12767 4646 12767 0 net17
rlabel metal1 4232 13498 4232 13498 0 net18
rlabel metal2 3266 14178 3266 14178 0 net19
rlabel metal2 11362 8160 11362 8160 0 net2
rlabel via3 4163 13804 4163 13804 0 net20
rlabel metal1 3358 14382 3358 14382 0 net21
rlabel metal1 2990 12954 2990 12954 0 net22
rlabel metal1 1426 7242 1426 7242 0 net23
rlabel metal1 10534 2414 10534 2414 0 net24
rlabel metal1 13018 11560 13018 11560 0 net3
rlabel via3 11293 13940 11293 13940 0 net4
rlabel metal2 13110 5032 13110 5032 0 net5
rlabel metal1 2392 2482 2392 2482 0 net6
rlabel metal2 2346 3706 2346 3706 0 net7
rlabel metal1 3588 3910 3588 3910 0 net8
rlabel metal1 4600 2414 4600 2414 0 net9
rlabel metal1 9016 14586 9016 14586 0 result[0]
rlabel metal1 7958 14586 7958 14586 0 result[1]
rlabel metal1 6992 14586 6992 14586 0 result[2]
rlabel metal1 5980 14586 5980 14586 0 result[3]
rlabel metal1 4968 14586 4968 14586 0 result[4]
rlabel metal1 3956 14586 3956 14586 0 result[5]
rlabel metal1 2944 14586 2944 14586 0 result[6]
rlabel metal1 1886 14586 1886 14586 0 result[7]
rlabel metal1 1150 14586 1150 14586 0 result_ready
rlabel metal1 13156 14382 13156 14382 0 rst
rlabel metal2 10442 1520 10442 1520 0 thresh_sel
rlabel metal1 10028 2414 10028 2414 0 use_ext_thresh
rlabel metal1 11040 14382 11040 14382 0 user_enable
rlabel metal1 13524 3706 13524 3706 0 wowa_digital.adc.comparator.compres.ffsync.stage0
rlabel metal1 6854 8942 6854 8942 0 wowa_digital.adc.comparator.compres.ffsync.stage1
rlabel metal1 10626 8466 10626 8466 0 wowa_digital.adc.internalCounter\[0\]
rlabel metal1 9522 9588 9522 9588 0 wowa_digital.adc.internalCounter\[1\]
rlabel metal1 8326 11730 8326 11730 0 wowa_digital.adc.internalCounter\[2\]
rlabel metal1 11546 13226 11546 13226 0 wowa_digital.adc.internalCounter\[3\]
rlabel metal1 9338 11662 9338 11662 0 wowa_digital.adc.internalCounter\[4\]
rlabel metal1 7974 13294 7974 13294 0 wowa_digital.adc.internalCounter\[5\]
rlabel metal1 8786 4556 8786 4556 0 wowa_digital.adc.state\[0\]
rlabel metal1 8050 6800 8050 6800 0 wowa_digital.adc.state\[1\]
rlabel metal1 11500 6766 11500 6766 0 wowa_digital.adc.state\[2\]
rlabel metal1 7314 6970 7314 6970 0 wowa_digital.adc.state\[3\]
rlabel metal1 9384 2414 9384 2414 0 wowa_digital.adc.syncroCount\[0\]
rlabel metal1 9384 2346 9384 2346 0 wowa_digital.adc.syncroCount\[1\]
<< properties >>
string FIXED_BBOX 0 0 15020 17164
<< end >>
