magic
tech sky130A
magscale 1 2
timestamp 1713335925
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 98 157 820 203
rect 1 21 820 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 188 47 218 177
rect 272 47 302 177
rect 460 47 490 177
rect 544 47 574 177
rect 628 47 658 177
rect 712 47 742 177
<< scpmoshvt >>
rect 79 413 109 497
rect 188 297 218 497
rect 272 297 302 497
rect 356 297 386 497
rect 440 297 470 497
rect 628 297 658 497
rect 712 297 742 497
<< ndiff >>
rect 124 161 188 177
rect 124 131 132 161
rect 27 101 79 131
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 127 132 131
rect 166 127 188 161
rect 109 93 188 127
rect 109 59 132 93
rect 166 59 188 93
rect 109 47 188 59
rect 218 161 272 177
rect 218 127 228 161
rect 262 127 272 161
rect 218 93 272 127
rect 218 59 228 93
rect 262 59 272 93
rect 218 47 272 59
rect 302 93 354 177
rect 302 59 312 93
rect 346 59 354 93
rect 302 47 354 59
rect 408 93 460 177
rect 408 59 416 93
rect 450 59 460 93
rect 408 47 460 59
rect 490 161 544 177
rect 490 127 500 161
rect 534 127 544 161
rect 490 47 544 127
rect 574 161 628 177
rect 574 127 584 161
rect 618 127 628 161
rect 574 93 628 127
rect 574 59 584 93
rect 618 59 628 93
rect 574 47 628 59
rect 658 169 712 177
rect 658 135 668 169
rect 702 135 712 169
rect 658 47 712 135
rect 742 93 794 177
rect 742 59 752 93
rect 786 59 794 93
rect 742 47 794 59
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 485 188 497
rect 109 451 132 485
rect 166 451 188 485
rect 109 417 188 451
rect 109 413 132 417
rect 124 383 132 413
rect 166 383 188 417
rect 124 297 188 383
rect 218 485 272 497
rect 218 451 228 485
rect 262 451 272 485
rect 218 417 272 451
rect 218 383 228 417
rect 262 383 272 417
rect 218 297 272 383
rect 302 485 356 497
rect 302 451 312 485
rect 346 451 356 485
rect 302 297 356 451
rect 386 485 440 497
rect 386 451 396 485
rect 430 451 440 485
rect 386 417 440 451
rect 386 383 396 417
rect 430 383 440 417
rect 386 297 440 383
rect 470 485 522 497
rect 470 451 480 485
rect 514 451 522 485
rect 470 297 522 451
rect 576 485 628 497
rect 576 451 584 485
rect 618 451 628 485
rect 576 297 628 451
rect 658 477 712 497
rect 658 443 668 477
rect 702 443 712 477
rect 658 409 712 443
rect 658 375 668 409
rect 702 375 712 409
rect 658 297 712 375
rect 742 485 794 497
rect 742 451 752 485
rect 786 451 794 485
rect 742 297 794 451
<< ndiffc >>
rect 35 67 69 101
rect 132 127 166 161
rect 132 59 166 93
rect 228 127 262 161
rect 228 59 262 93
rect 312 59 346 93
rect 416 59 450 93
rect 500 127 534 161
rect 584 127 618 161
rect 584 59 618 93
rect 668 135 702 169
rect 752 59 786 93
<< pdiffc >>
rect 35 443 69 477
rect 132 451 166 485
rect 132 383 166 417
rect 228 451 262 485
rect 228 383 262 417
rect 312 451 346 485
rect 396 451 430 485
rect 396 383 430 417
rect 480 451 514 485
rect 584 451 618 485
rect 668 443 702 477
rect 668 375 702 409
rect 752 451 786 485
<< poly >>
rect 79 497 109 523
rect 188 497 218 523
rect 272 497 302 523
rect 356 497 386 523
rect 440 497 470 523
rect 628 497 658 523
rect 712 497 742 523
rect 79 265 109 413
rect 79 249 146 265
rect 79 215 102 249
rect 136 215 146 249
rect 79 199 146 215
rect 188 259 218 297
rect 272 259 302 297
rect 188 249 302 259
rect 188 215 228 249
rect 262 215 302 249
rect 188 205 302 215
rect 356 259 386 297
rect 440 259 470 297
rect 628 259 658 297
rect 712 259 742 297
rect 356 249 574 259
rect 356 215 406 249
rect 440 215 478 249
rect 512 215 574 249
rect 356 205 574 215
rect 79 131 109 199
rect 188 177 218 205
rect 272 177 302 205
rect 460 177 490 205
rect 544 177 574 205
rect 628 249 742 259
rect 628 215 680 249
rect 714 215 742 249
rect 628 205 742 215
rect 628 177 658 205
rect 712 177 742 205
rect 79 21 109 47
rect 188 21 218 47
rect 272 21 302 47
rect 460 21 490 47
rect 544 21 574 47
rect 628 21 658 47
rect 712 21 742 47
<< polycont >>
rect 102 215 136 249
rect 228 215 262 249
rect 406 215 440 249
rect 478 215 512 249
rect 680 215 714 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 477 82 493
rect 18 443 35 477
rect 69 443 82 477
rect 18 413 82 443
rect 116 485 178 527
rect 116 451 132 485
rect 166 451 178 485
rect 116 417 178 451
rect 18 323 52 413
rect 116 383 132 417
rect 166 383 178 417
rect 116 367 178 383
rect 212 485 278 493
rect 212 451 228 485
rect 262 451 278 485
rect 212 417 278 451
rect 312 485 346 527
rect 312 435 346 451
rect 380 485 446 493
rect 380 451 396 485
rect 430 451 446 485
rect 212 383 228 417
rect 262 401 278 417
rect 380 417 446 451
rect 480 485 530 527
rect 514 451 530 485
rect 480 435 530 451
rect 568 485 618 527
rect 568 451 584 485
rect 568 435 618 451
rect 652 477 702 493
rect 652 443 668 477
rect 380 401 396 417
rect 262 383 396 401
rect 430 391 446 417
rect 652 409 702 443
rect 752 485 810 527
rect 786 451 810 485
rect 752 435 810 451
rect 652 391 668 409
rect 430 383 668 391
rect 212 375 668 383
rect 702 375 810 401
rect 212 357 810 375
rect 18 289 730 323
rect 18 131 52 289
rect 86 249 156 255
rect 86 215 102 249
rect 136 215 156 249
rect 212 249 348 255
rect 212 215 228 249
rect 262 215 348 249
rect 390 249 628 255
rect 390 215 406 249
rect 440 215 478 249
rect 512 215 628 249
rect 664 249 730 289
rect 664 215 680 249
rect 714 215 730 249
rect 770 181 810 357
rect 116 161 178 181
rect 18 101 82 131
rect 18 67 35 101
rect 69 67 82 101
rect 18 51 82 67
rect 116 127 132 161
rect 166 127 178 161
rect 116 93 178 127
rect 116 59 132 93
rect 166 59 178 93
rect 116 17 178 59
rect 212 161 550 181
rect 212 127 228 161
rect 262 143 500 161
rect 262 127 278 143
rect 400 127 500 143
rect 534 127 550 161
rect 584 161 618 181
rect 652 169 810 181
rect 652 135 668 169
rect 702 135 810 169
rect 652 127 810 135
rect 212 93 278 127
rect 212 59 228 93
rect 262 59 278 93
rect 212 51 278 59
rect 312 93 362 109
rect 584 93 618 127
rect 346 59 362 93
rect 312 17 362 59
rect 400 59 416 93
rect 450 59 584 93
rect 618 59 752 93
rect 786 59 810 93
rect 400 51 810 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 C
port 7 nsew
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A_N
port 6 nsew
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 B
port 8 nsew
flabel locali s 770 289 804 323 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel locali s 415 238 415 238 0 FreeSans 200 0 0 0 B
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 nand3b_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 216752
string GDS_FILE wowa_digital_ol.gds
string GDS_START 209804
string path 0.000 0.000 4.140 0.000 
<< end >>
