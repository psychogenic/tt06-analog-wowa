magic
tech sky130A
magscale 1 2
timestamp 1713150084
<< metal4 >>
rect -1849 8339 1849 8380
rect -1849 5261 1593 8339
rect 1829 5261 1849 8339
rect -1849 5220 1849 5261
rect -1849 4939 1849 4980
rect -1849 1861 1593 4939
rect 1829 1861 1849 4939
rect -1849 1820 1849 1861
rect -1849 1539 1849 1580
rect -1849 -1539 1593 1539
rect 1829 -1539 1849 1539
rect -1849 -1580 1849 -1539
rect -1849 -1861 1849 -1820
rect -1849 -4939 1593 -1861
rect 1829 -4939 1849 -1861
rect -1849 -4980 1849 -4939
rect -1849 -5261 1849 -5220
rect -1849 -8339 1593 -5261
rect 1829 -8339 1849 -5261
rect -1849 -8380 1849 -8339
<< via4 >>
rect 1593 5261 1829 8339
rect 1593 1861 1829 4939
rect 1593 -1539 1829 1539
rect 1593 -4939 1829 -1861
rect 1593 -8339 1829 -5261
<< mimcap2 >>
rect -1769 8260 1231 8300
rect -1769 5340 -1729 8260
rect 1191 5340 1231 8260
rect -1769 5300 1231 5340
rect -1769 4860 1231 4900
rect -1769 1940 -1729 4860
rect 1191 1940 1231 4860
rect -1769 1900 1231 1940
rect -1769 1460 1231 1500
rect -1769 -1460 -1729 1460
rect 1191 -1460 1231 1460
rect -1769 -1500 1231 -1460
rect -1769 -1940 1231 -1900
rect -1769 -4860 -1729 -1940
rect 1191 -4860 1231 -1940
rect -1769 -4900 1231 -4860
rect -1769 -5340 1231 -5300
rect -1769 -8260 -1729 -5340
rect 1191 -8260 1231 -5340
rect -1769 -8300 1231 -8260
<< mimcap2contact >>
rect -1729 5340 1191 8260
rect -1729 1940 1191 4860
rect -1729 -1460 1191 1460
rect -1729 -4860 1191 -1940
rect -1729 -8260 1191 -5340
<< metal5 >>
rect -429 8284 -109 8500
rect 1551 8339 1871 8500
rect -1753 8260 1215 8284
rect -1753 5340 -1729 8260
rect 1191 5340 1215 8260
rect -1753 5316 1215 5340
rect -429 4884 -109 5316
rect 1551 5261 1593 8339
rect 1829 5261 1871 8339
rect 1551 4939 1871 5261
rect -1753 4860 1215 4884
rect -1753 1940 -1729 4860
rect 1191 1940 1215 4860
rect -1753 1916 1215 1940
rect -429 1484 -109 1916
rect 1551 1861 1593 4939
rect 1829 1861 1871 4939
rect 1551 1539 1871 1861
rect -1753 1460 1215 1484
rect -1753 -1460 -1729 1460
rect 1191 -1460 1215 1460
rect -1753 -1484 1215 -1460
rect -429 -1916 -109 -1484
rect 1551 -1539 1593 1539
rect 1829 -1539 1871 1539
rect 1551 -1861 1871 -1539
rect -1753 -1940 1215 -1916
rect -1753 -4860 -1729 -1940
rect 1191 -4860 1215 -1940
rect -1753 -4884 1215 -4860
rect -429 -5316 -109 -4884
rect 1551 -4939 1593 -1861
rect 1829 -4939 1871 -1861
rect 1551 -5261 1871 -4939
rect -1753 -5340 1215 -5316
rect -1753 -8260 -1729 -5340
rect 1191 -8260 1215 -5340
rect -1753 -8284 1215 -8260
rect -429 -8500 -109 -8284
rect 1551 -8339 1593 -5261
rect 1829 -8339 1871 -5261
rect 1551 -8500 1871 -8339
<< properties >>
string FIXED_BBOX -1849 5220 1311 8380
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 15.0 l 15.0 val 461.4 carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
