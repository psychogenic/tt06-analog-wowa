magic
tech sky130A
magscale 1 2
timestamp 1713123902
<< error_p >>
rect -29 272 29 278
rect -29 238 -17 272
rect -29 232 29 238
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect -29 -278 29 -272
<< pwell >>
rect -216 -410 216 410
<< nmos >>
rect -20 -200 20 200
<< ndiff >>
rect -78 188 -20 200
rect -78 -188 -66 188
rect -32 -188 -20 188
rect -78 -200 -20 -188
rect 20 188 78 200
rect 20 -188 32 188
rect 66 -188 78 188
rect 20 -200 78 -188
<< ndiffc >>
rect -66 -188 -32 188
rect 32 -188 66 188
<< psubdiff >>
rect -180 340 -84 374
rect 84 340 180 374
rect -180 278 -146 340
rect 146 278 180 340
rect -180 -340 -146 -278
rect 146 -340 180 -278
rect -180 -374 -84 -340
rect 84 -374 180 -340
<< psubdiffcont >>
rect -84 340 84 374
rect -180 -278 -146 278
rect 146 -278 180 278
rect -84 -374 84 -340
<< poly >>
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect -20 200 20 222
rect -20 -222 20 -200
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -180 340 -84 374
rect 84 340 180 374
rect -180 278 -146 340
rect 146 278 180 340
rect -33 238 -17 272
rect 17 238 33 272
rect -66 188 -32 204
rect -66 -204 -32 -188
rect 32 188 66 204
rect 32 -204 66 -188
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -180 -340 -146 -278
rect 146 -340 180 -278
rect -180 -374 -84 -340
rect 84 -374 180 -340
<< viali >>
rect -17 238 17 272
rect -66 -188 -32 188
rect 32 -188 66 188
rect -17 -272 17 -238
<< metal1 >>
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect -72 188 -26 200
rect -72 -188 -66 188
rect -32 -188 -26 188
rect -72 -200 -26 -188
rect 26 188 72 200
rect 26 -188 32 188
rect 66 -188 72 188
rect 26 -200 72 -188
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
<< properties >>
string FIXED_BBOX -163 -357 163 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
