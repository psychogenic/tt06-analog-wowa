** sch_path: /home/ttuser/wowa/xschem/wowa_analog.sch
.subckt wowa_analog b0 b1 b2 b3 b4 b5 b6 b7 EN_N CAL INPUT EXTTHRESH USEEXT VCC VSS COMPOUT
*.PININFO b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I EN_N:I CAL:I INPUT:I EXTTHRESH:I USEEXT:I VCC:I
*+ VSS:I COMPOUT:O
x1 VCC VSS INPUT THRESH COMPOUT CAL EN_N calibrated_comparator
x2 b0 b1 b2 b3 b4 b5 b6 b7 INTTHRESH VSS VSS r2r
x3 VCC VSS USEEXT EXTTHRESH THRESH INTTHRESH onehot2mux
.ends

* expanding   symbol:  /home/ttuser/wowa/xschem/calibrated_comparator.sym # of pins=7
** sym_path: /home/ttuser/wowa/xschem/calibrated_comparator.sym
** sch_path: /home/ttuser/wowa/xschem/calibrated_comparator.sch
.subckt calibrated_comparator VCC VSS INPUT THRESHV RESULT CALIB EN_N
*.PININFO VCC:I VSS:I INPUT:I THRESHV:I CALIB:I RESULT:O EN_N:I
x1 VCC VSS EN_N ADJ RESULT INSIG THRESHV comparator_stefan
x2 VCC VSS CALIB ADJ RESULT analogswitch
x3 VCC VSS CALIB THRESHV INSIG INPUT onehot2mux
XC1 ADJ VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=4
.ends


* expanding   symbol:  /home/ttuser/wowa/tt06-analog-r2r-dac/xschem/r2r.sym # of pins=11
** sym_path: /home/ttuser/wowa/tt06-analog-r2r-dac/xschem/r2r.sym
** sch_path: /home/ttuser/wowa/tt06-analog-r2r-dac/xschem/r2r.sch
.subckt r2r b0 b1 b2 b3 b4 b5 b6 b7 out GND VSUBS
*.PININFO b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I out:O VSUBS:I GND:B
XR1 net1 b0 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR2 net2 b1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR3 net3 b2 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR4 net4 b3 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR5 net5 b4 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR6 net6 b5 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR7 net7 b6 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR8 out b7 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
XR9 net2 net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR10 net3 net2 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR11 net4 net3 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR12 net5 net4 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR13 net6 net5 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR14 net7 net6 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR15 out net7 VSUBS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XR16 GND net1 VSUBS sky130_fd_pr__res_high_po_0p35 L=40 mult=1 m=1
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/onehot2mux.sym # of pins=6
** sym_path: /home/ttuser/wowa/xschem/onehot2mux.sym
** sch_path: /home/ttuser/wowa/xschem/onehot2mux.sch
.subckt onehot2mux VCC VSS SEL IN1 OUT IN0
*.PININFO SEL:I IN0:I IN1:I OUT:O VCC:I VSS:I
x2 OUT IN1 SEL_N SEL VSS VCC passgate
x3 OUT IN0 SEL SEL_N VSS VCC passgate
x1 SEL SEL_N VCC VSS lvtnot
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/comparator_stefan.sym # of pins=7
** sym_path: /home/ttuser/wowa/xschem/comparator_stefan.sym
** sch_path: /home/ttuser/wowa/xschem/comparator_stefan.sch
.subckt comparator_stefan VCC VSS EN_N ADJ DIFFOUT PLUS MINUS
*.PININFO PLUS:I MINUS:I VCC:I VSS:I EN_N:I ADJ:I DIFFOUT:O
XM1 inhigh EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=2 nf=1 m=1
XM2 G1 MINUS inhigh VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 m=1
XM3 inhigh PLUS G2 VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 m=1
XM4 G2 G2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM5 VSS G1 G1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM6 pg2g G1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM7 mirhigh pg2g pg2g VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 m=1
XM8 DIFFOUT pg2g mirhigh VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 m=1
XM9 mirhigh EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 m=1
XM10 DIFFOUT G2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 m=1
XM11 DIFFOUT EN_N VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 p2p EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM13 G1 ADJ p2p VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM14 G1 ADJ n2n VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.5 nf=1 m=1
XM15 n2n VCC VSS VSS sky130_fd_pr__nfet_01v8_lvt L=8 W=0.5 nf=1 m=1
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/analogswitch.sym # of pins=5
** sym_path: /home/ttuser/wowa/xschem/analogswitch.sym
** sch_path: /home/ttuser/wowa/xschem/analogswitch.sch
.subckt analogswitch VCC VSS EN OUT IN
*.PININFO EN:I IN:I OUT:O VCC:I VSS:I
x2 OUT IN EN_N EN VSS VCC passgate
x1 EN EN_N VCC VSS lvtnot
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/wowa/xschem/passgate.sym
** sch_path: /home/ttuser/wowa/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.PININFO A:B Z:B GP:I GN:I VCCBPIN:I VSSBPIN:I
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8 L=0.2 W=2 nf=1 m=1
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/lvtnot.sym # of pins=4
** sym_path: /home/ttuser/wowa/xschem/lvtnot.sym
** sch_path: /home/ttuser/wowa/xschem/lvtnot.sch
.subckt lvtnot a y VCCPIN VSSPIN
*.PININFO y:O a:I VCCPIN:I VSSPIN:I
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 m=1
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
.ends

.end
