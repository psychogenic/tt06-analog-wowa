* NGSPICE file created from lvtnot_parax.ext - technology: sky130A

.subckt lvtnot_parax a y VCCPIN VSSPIN
X0 VCCPIN.t1 a.t0 y.t0 VCCPIN.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
X1 y.t1 a.t1 VSSPIN.t1 VSSPIN.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 a.n0 a.t1 193.226
R1 a.n0 a.t0 174.12
R2 a a.n0 1.188
R3 y.n0 y.t0 113.802
R4 y.n0 y.t1 83.8505
R5 y y.n0 0.20699
R6 VCCPIN.n8 VCCPIN.n2 1860
R7 VCCPIN.n6 VCCPIN.n5 1860
R8 VCCPIN.n5 VCCPIN.n4 561.481
R9 VCCPIN.n8 VCCPIN.n7 561.481
R10 VCCPIN.n9 VCCPIN.n1 198.4
R11 VCCPIN.n3 VCCPIN.n1 198.4
R12 VCCPIN.n3 VCCPIN.n0 175.391
R13 VCCPIN.n10 VCCPIN.n9 173.403
R14 VCCPIN.n11 VCCPIN.t1 113.645
R15 VCCPIN.n9 VCCPIN.n8 61.6672
R16 VCCPIN.n5 VCCPIN.n3 61.6672
R17 VCCPIN.n6 VCCPIN.n1 23.1255
R18 VCCPIN.n2 VCCPIN.n0 23.1255
R19 VCCPIN.n4 VCCPIN.n2 15.947
R20 VCCPIN.n7 VCCPIN.n6 15.947
R21 VCCPIN.n7 VCCPIN.t0 6.98177
R22 VCCPIN.n4 VCCPIN.t0 6.98177
R23 VCCPIN.n11 VCCPIN.n10 1.8605
R24 VCCPIN.n10 VCCPIN.n0 1.0245
R25 VCCPIN.n12 VCCPIN 0.124875
R26 VCCPIN VCCPIN.n12 0.109601
R27 VCCPIN.n12 VCCPIN.n11 0.107956
R28 VSSPIN.n5 VSSPIN.n3 2306.06
R29 VSSPIN.n8 VSSPIN.n2 2306.06
R30 VSSPIN.n6 VSSPIN.n2 1183.39
R31 VSSPIN.n7 VSSPIN.n3 1183.39
R32 VSSPIN.n2 VSSPIN.n1 292.5
R33 VSSPIN.n3 VSSPIN.n0 292.5
R34 VSSPIN.n4 VSSPIN.n1 149.835
R35 VSSPIN.n4 VSSPIN.n0 149.835
R36 VSSPIN.n9 VSSPIN.n1 126.947
R37 VSSPIN.n10 VSSPIN.n0 124.462
R38 VSSPIN.n5 VSSPIN.n4 117.001
R39 VSSPIN.n9 VSSPIN.n8 117.001
R40 VSSPIN.n11 VSSPIN.t1 83.7278
R41 VSSPIN.n7 VSSPIN.t0 60.0412
R42 VSSPIN.t0 VSSPIN.n6 60.0412
R43 VSSPIN.n6 VSSPIN.n5 54.2104
R44 VSSPIN.n8 VSSPIN.n7 54.2104
R45 VSSPIN.n11 VSSPIN.n10 1.86348
R46 VSSPIN.n10 VSSPIN.n9 1.2805
R47 VSSPIN VSSPIN.n11 0.244548
C0 y VCCPIN 0.488784f
C1 y a 0.532131f
C2 a VCCPIN 0.819808f
C3 y VSSPIN 0.541674f
C4 a VSSPIN 1.46791f
C5 VCCPIN VSSPIN 1.99105f
.ends

