magic
tech sky130A
magscale 1 2
timestamp 1713420955
<< locali >>
rect 2410 1290 3050 1310
rect 2410 1200 2500 1290
rect 2980 1200 3050 1290
rect 2410 1150 3050 1200
rect 2410 1110 2590 1150
rect 2840 1110 3050 1150
rect 2880 1050 3050 1110
rect 2900 970 3050 1050
rect 2880 940 3050 970
rect 2460 -440 2560 -230
rect 2870 -290 2970 -230
rect 2870 -300 3110 -290
rect 2900 -380 3110 -300
rect 2200 -470 2590 -440
rect 2870 -440 3110 -380
rect 2840 -470 3110 -440
rect 2200 -540 3110 -470
rect 2200 -650 2330 -540
rect 3050 -650 3110 -540
rect 2200 -700 3110 -650
<< viali >>
rect 2500 1200 2980 1290
rect 2590 1110 2840 1150
rect 2860 970 2900 1050
rect 2860 -380 2900 -300
rect 2590 -470 2840 -430
rect 2330 -650 3050 -540
<< metal1 >>
rect 2200 1290 3110 1400
rect 2200 1200 2500 1290
rect 2980 1200 3110 1290
rect 2200 1150 3110 1200
rect 2200 1130 2590 1150
rect 2500 1110 2590 1130
rect 2840 1110 3110 1150
rect 2500 1100 3110 1110
rect 2200 1047 2400 1100
rect 2840 1050 3110 1100
rect 2200 954 2373 1047
rect 2466 954 2472 1047
rect 2680 990 2690 1050
rect 2750 990 2760 1050
rect 2840 970 2860 1050
rect 2900 970 3110 1050
rect 2200 900 2400 954
rect 2840 940 3110 970
rect 2490 810 2690 880
rect 2330 570 2690 810
rect 2750 810 2950 880
rect 2750 570 3110 810
rect 2330 500 2550 570
rect 2200 300 2550 500
rect 2680 460 2690 520
rect 2750 460 2760 520
rect 2890 500 3110 570
rect 2330 100 2550 300
rect 2890 300 3200 500
rect 2670 140 2680 210
rect 2760 140 2770 210
rect 2890 100 3110 300
rect 2330 -130 2690 100
rect 2200 -301 2400 -200
rect 2490 -210 2690 -130
rect 2740 -130 3110 100
rect 2740 -210 2940 -130
rect 2840 -300 3110 -290
rect 2200 -307 2487 -301
rect 2200 -400 2394 -307
rect 2670 -390 2680 -320
rect 2760 -390 2770 -320
rect 2840 -380 2860 -300
rect 2900 -380 3110 -300
rect 2394 -406 2487 -400
rect 2840 -420 3110 -380
rect 2540 -430 3110 -420
rect 2540 -440 2590 -430
rect 2200 -470 2590 -440
rect 2840 -470 3110 -430
rect 2200 -540 3110 -470
rect 2200 -650 2330 -540
rect 3050 -650 3110 -540
rect 2200 -700 3110 -650
<< via1 >>
rect 2373 954 2466 1047
rect 2690 990 2750 1050
rect 2690 460 2750 520
rect 2680 140 2760 210
rect 2394 -400 2487 -307
rect 2680 -390 2760 -320
<< metal2 >>
rect 2373 1047 2466 1053
rect 2680 1050 2760 1060
rect 2680 1047 2690 1050
rect 2466 990 2690 1047
rect 2750 1047 2760 1050
rect 2750 990 2766 1047
rect 2466 954 2766 990
rect 2373 948 2466 954
rect 2673 520 2766 954
rect 2673 460 2690 520
rect 2750 460 2766 520
rect 2673 454 2766 460
rect 2690 450 2750 454
rect 2673 210 2766 226
rect 2673 140 2680 210
rect 2760 140 2766 210
rect 2673 -307 2766 140
rect 2388 -400 2394 -307
rect 2487 -320 2766 -307
rect 2487 -390 2680 -320
rect 2760 -390 2766 -320
rect 2487 -400 2766 -390
use sky130_fd_pr__nfet_01v8_Q7AWK3  XM1
timestamp 1713123902
transform 1 0 2716 0 1 -90
box -216 -410 216 410
use sky130_fd_pr__pfet_01v8_SKB8XJ  XM2
timestamp 1713123902
transform -1 0 2716 0 -1 759
box -216 -419 216 419
<< labels >>
flabel metal1 2200 -400 2400 -200 0 FreeSans 1280 0 0 0 GN
port 3 nsew
flabel metal1 3000 300 3200 500 0 FreeSans 1280 0 0 0 Z
port 1 nsew
flabel metal1 2200 300 2400 500 0 FreeSans 1280 0 0 0 A
port 0 nsew
flabel metal1 2200 900 2400 1100 0 FreeSans 1280 0 0 0 GP
port 2 nsew
flabel metal1 2600 -700 2800 -500 0 FreeSans 1280 0 0 0 VSSBPIN
port 5 nsew
flabel metal1 2600 1200 2800 1400 0 FreeSans 1280 0 0 0 VCCBPIN
port 4 nsew
<< end >>
