** sch_path: /home/ttuser/wowa/xschem/analogswitch.sch
.subckt analogswitch EN IN OUT VCC VSS
*.PININFO EN:I IN:I OUT:O VCC:I VSS:I
x2 OUT IN EN_N EN VSS VCC passgate
x1 EN EN_N VCC VSS lvtnot
.ends

* expanding   symbol:  /home/ttuser/wowa/xschem/passgate.sym # of pins=6
** sym_path: /home/ttuser/wowa/xschem/passgate.sym
** sch_path: /home/ttuser/wowa/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.PININFO A:B Z:B GP:I GN:I VCCBPIN:I VSSBPIN:I
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8 L=0.2 W=2 nf=1 m=1
.ends


* expanding   symbol:  /home/ttuser/wowa/xschem/lvtnot.sym # of pins=4
** sym_path: /home/ttuser/wowa/xschem/lvtnot.sym
** sch_path: /home/ttuser/wowa/xschem/lvtnot.sch
.subckt lvtnot a y VCCPIN VSSPIN
*.PININFO y:O a:I VCCPIN:I VSSPIN:I
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 m=1
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
.ends

.end
