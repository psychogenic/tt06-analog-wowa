** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/tb_calibrated_comparator_eyediag.sch
**.subckt tb_calibrated_comparator_eyediag
x1 VCC VSS INPUT THRESHV RESULT CALIB EN_N calibrated_comparator
x2 VCC VSS INPUT THRESHV RESULT_PARAX CALIB EN_N calibrated_comparator
XR1 INPUT_A INPUT net1 sky130_fd_pr__res_xhigh_po_1p41 L=40 mult=1 m=1
XR2 INPUT_B INPUT net2 sky130_fd_pr__res_xhigh_po_1p41 L=40 mult=1 m=1
VINPULSE INPUT_B VSS pulse VLOW VHIGH 1u 5n 5n PULSEWIDTH PULSEPER
VTH THRESHV VSS dc 0.6
**** begin user architecture code

.param mc_mm_switch=1
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



** this experimental option enables mos model bin
** selection based on W/NF instead of W
.option chgtol=4e-16 method=gear

.param VCCGAUSS = agauss(1.8, 0.05, 1)
.param VCC = 'VCCGAUSS'
** use following line to remove VCC variations
* .param VCC = 1.8
.param VDLGAUSS = agauss(0.9, 0.23, 1)
.param VDL = VDLGAUSS
** use following line to remove input common mode variations
* .param VDL =  1.4
.param TEMPGAUSS = agauss(40, 30, 1)
.option temp = 'TEMPGAUSS'
** use following line to remove temperature variations
* .option temp = 25
.param DELTA = 0.002


* VLOW VHIGH 900n 1n 1n PULSEWIDTH PULSEPER


* our calibration stage/setup
.include stimuli_tb_calibrated_comparator_eyediag.cir

.param VLOW = -0.2
.param VHIGH =2.2
.param PULSEWIDTH = 100n
.param PULSEPER = 200n


.control
  setseed  8
  reset
  let run = 1
  let pw = 50n
  let pp = 100n
  let vthresh = 0.01
  save all
  op
  write tb_calibrated_comparator_eyediag.raw
  reset
  set appendwrite
  dowhile vthresh <= 1.6

   alter VTH vthresh
   dowhile run < = 3
    save all
    let pw = pw * 2
    let pp = pw * 2
    * alter VINPULSE PW = pw
    * alter VINPULSE PER = pp
    tran 1n 3200n uic
    write tb_calibrated_comparator_eyediag.raw
    let run = run + 1
    reset
   end
   let vthresh = vthresh + 0.05
  end
  quit 0
.endc


**** end user architecture code
**.ends

* expanding   symbol:  calibrated_comparator.sym # of pins=7
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/calibrated_comparator.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/calibrated_comparator.sch
.subckt calibrated_comparator VCC VSS INPUT THRESHV RESULT CALIB EN_N
*.ipin VCC
*.ipin VSS
*.ipin INPUT
*.ipin THRESHV
*.ipin CALIB
*.opin RESULT
*.ipin EN_N
x1 VCC VSS EN_N ADJ RESULT INSIG THRESHV comparator_stefan
x2 VCC VSS CALIB ADJ RESULT analogswitch
x3 VCC VSS CALIB THRESHV INSIG INPUT onehot2mux
XC1 ADJ VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
.ends


* expanding   symbol:  comparator_stefan.sym # of pins=7
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/comparator_stefan.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/comparator_stefan.sch
.subckt comparator_stefan VCC VSS EN_N ADJ DIFFOUT PLUS MINUS
*.ipin PLUS
*.ipin MINUS
*.ipin VCC
*.ipin VSS
*.ipin EN_N
*.ipin ADJ
*.opin DIFFOUT
XM1 inhigh EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 G1 MINUS inhigh VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 inhigh PLUS G2 VCC sky130_fd_pr__pfet_01v8_lvt L=2 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 G2 G2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 VSS G1 G1 VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 pg2g G1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 mirhigh pg2g pg2g VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 DIFFOUT pg2g mirhigh VCC sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 mirhigh EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 DIFFOUT G2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 DIFFOUT EN_N VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 p2p EN_N VCC VCC sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 G1 ADJ p2p VCC sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 G1 ADJ n2n VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM15 n2n VCC VSS VSS sky130_fd_pr__nfet_01v8_lvt L=8 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  analogswitch.sym # of pins=5
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/analogswitch.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/analogswitch.sch
.subckt analogswitch VCC VSS EN OUT IN
*.ipin EN
*.ipin IN
*.opin OUT
*.ipin VCC
*.ipin VSS
x2 OUT IN EN_N EN VSS VCC passgate
x1 EN EN_N VCC VSS lvtnot
.ends


* expanding   symbol:  onehot2mux.sym # of pins=6
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/onehot2mux.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/onehot2mux.sch
.subckt onehot2mux VCC VSS SEL IN1 OUT IN0
*.ipin SEL
*.ipin IN0
*.ipin IN1
*.opin OUT
*.ipin VCC
*.ipin VSS
x2 OUT IN1 SEL_N SEL VSS VCC passgate
x3 OUT IN0 SEL SEL_N VSS VCC passgate
x1 SEL SEL_N VCC VSS lvtnot
.ends


* expanding   symbol:  passgate.sym # of pins=6
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/passgate.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/passgate.sch
.subckt passgate Z A GP GN VSSBPIN VCCBPIN
*.iopin A
*.iopin Z
*.ipin GP
*.ipin GN
*.ipin VCCBPIN
*.ipin VSSBPIN
XM1 Z GN A VSSBPIN sky130_fd_pr__nfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z GP A VCCBPIN sky130_fd_pr__pfet_01v8 L=0.2 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  lvtnot.sym # of pins=4
** sym_path: /home/ttuser/work/tt06-analog-wowa/xschem/lvtnot.sym
** sch_path: /home/ttuser/work/tt06-analog-wowa/xschem/lvtnot.sch
.subckt lvtnot a y VCCPIN VSSPIN
*.opin y
*.ipin a
*.ipin VCCPIN
*.ipin VSSPIN
XM2 y a VCCPIN VCCPIN sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 y a VSSPIN VSSPIN sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
