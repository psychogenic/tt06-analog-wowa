magic
tech sky130A
magscale 1 2
timestamp 1713301548
<< metal1 >>
rect 23560 19159 29606 19206
rect 23560 18961 23631 19159
rect 23829 18961 29606 19159
rect 23560 18873 29606 18961
rect 6094 17890 6100 18450
rect 6660 17890 7300 18450
rect 7658 18442 7862 18448
rect 7538 18238 7658 18442
rect 8237 18303 8243 18497
rect 8437 18303 8443 18497
rect 8828 18295 8834 18506
rect 9045 18295 9051 18506
rect 9436 18302 9442 18498
rect 9638 18302 9644 18498
rect 9896 18296 10096 18504
rect 10304 18296 10310 18504
rect 10707 18493 10893 18499
rect 10507 18307 10707 18493
rect 11333 18323 11339 18477
rect 11493 18323 11499 18477
rect 11929 18335 11935 18465
rect 12065 18335 12071 18465
rect 10707 18301 10893 18307
rect 12566 18282 12572 18498
rect 12788 18282 12794 18498
rect 7658 18232 7862 18238
rect 12572 17942 12788 18282
rect 14018 18274 14024 18466
rect 14216 18274 14222 18466
rect 21622 18289 21628 18492
rect 21831 18289 21837 18492
rect 14024 17944 14216 18274
rect 21628 17929 21831 18289
rect 23586 18260 23867 18873
rect 14754 17440 14760 17840
rect 15160 17440 15166 17840
rect 22414 17440 22420 17840
rect 22820 17440 22826 17840
rect 14760 16640 15160 17440
rect 22420 17080 22820 17440
rect 15850 12680 15860 12860
rect 16300 12680 16310 12860
rect 21150 12660 21160 12920
rect 21480 12660 21490 12920
rect 16950 9320 16960 9420
rect 18740 9320 18750 9420
rect 21770 9260 21780 9360
rect 22360 9260 22370 9360
rect 25671 8069 26089 8075
rect 25671 7645 26089 7651
rect 25744 6924 27120 7277
rect 14010 4100 14020 4400
rect 14240 4100 14250 4400
rect 15360 4060 15700 4540
rect 12030 3620 12040 3860
rect 12300 3620 12310 3860
rect 6450 3060 6460 3200
rect 6980 3060 6990 3200
rect 15910 3116 16202 3286
rect 15881 2916 16232 3116
rect 21530 3000 21540 3260
rect 21900 3000 21910 3260
rect 25390 3000 25400 3280
rect 25860 3000 25870 3280
rect 15881 2565 16232 2655
rect 26752 940 27105 6924
rect 26752 700 26800 940
rect 27060 700 27105 940
rect 26752 644 27105 700
rect 29273 987 29606 18873
rect 29273 983 31366 987
rect 29273 960 31583 983
rect 29273 680 31280 960
rect 31540 680 31583 960
rect 29273 657 31583 680
rect 29273 654 31366 657
<< via1 >>
rect 23631 18961 23829 19159
rect 6100 17890 6660 18450
rect 7658 18238 7862 18442
rect 8243 18303 8437 18497
rect 8834 18295 9045 18506
rect 9442 18302 9638 18498
rect 10096 18296 10304 18504
rect 10707 18307 10893 18493
rect 11339 18323 11493 18477
rect 11935 18335 12065 18465
rect 12572 18282 12788 18498
rect 14024 18274 14216 18466
rect 21628 18289 21831 18492
rect 14760 17440 15160 17840
rect 22420 17440 22820 17840
rect 15860 12680 16300 12860
rect 21160 12660 21480 12920
rect 16960 9320 18740 9420
rect 21780 9260 22360 9360
rect 25671 7651 26089 8069
rect 14020 4100 14240 4400
rect 12040 3620 12300 3860
rect 6460 3060 6980 3200
rect 21540 3000 21900 3260
rect 25400 3000 25860 3280
rect 15881 2655 16232 2916
rect 26800 700 27060 940
rect 31280 680 31540 960
<< metal2 >>
rect 5211 44900 12558 44981
rect 5211 44898 9620 44900
rect 9780 44898 12558 44900
rect 12641 44898 12650 44981
rect 4191 43569 4290 43578
rect 4191 41451 4290 43470
rect 5211 41539 5294 44898
rect 9621 44794 9704 44800
rect 6230 44725 13305 44794
rect 13374 44725 13383 44794
rect 6230 41526 6299 44725
rect 9621 44719 9704 44725
rect 7241 44584 14044 44655
rect 14115 44584 14124 44655
rect 7241 41505 7312 44584
rect 8253 44445 14765 44515
rect 14835 44445 14844 44515
rect 8253 41505 8323 44445
rect 9259 44278 15498 44361
rect 15581 44278 15590 44361
rect 9259 41499 9342 44278
rect 16236 44164 16324 44173
rect 10268 44076 16236 44164
rect 10268 41496 10356 44076
rect 16236 44067 16324 44076
rect 11279 43957 17062 43962
rect 11279 43884 16984 43957
rect 17057 43884 17066 43957
rect 11279 43879 17062 43884
rect 11279 41519 11362 43879
rect 17724 43815 17795 43824
rect 12301 43744 17724 43775
rect 12301 43704 17795 43744
rect 12301 41505 12372 43704
rect 28016 43683 28103 43692
rect 28016 43583 28103 43596
rect 13305 43496 28103 43583
rect 13305 41477 13392 43496
rect 28733 43407 28827 43416
rect 14313 43313 28733 43327
rect 14313 43233 28827 43313
rect 14313 41453 14407 43233
rect 29497 42903 29583 42912
rect 15329 42817 29497 42903
rect 15329 41457 15415 42817
rect 29497 42808 29583 42817
rect 16330 42093 27060 42095
rect 16330 42082 27377 42093
rect 16330 41998 27282 42082
rect 27366 41998 27377 42082
rect 16330 41988 27377 41998
rect 16330 41986 27060 41988
rect 16345 41481 16423 41986
rect 30953 41747 31047 41756
rect 30953 41627 31047 41653
rect 17349 41533 31047 41627
rect 4138 21362 4342 24882
rect 5339 22097 5533 24817
rect 6527 22746 6738 24806
rect 7730 23358 7926 24858
rect 8920 24104 9128 24904
rect 8920 23896 9704 24104
rect 7730 23162 9078 23358
rect 6527 22535 8445 22746
rect 5339 21903 7797 22097
rect 4138 21158 7102 21362
rect 6100 18450 6660 18456
rect 1191 17890 1200 18450
rect 1760 17890 6100 18450
rect 6898 18442 7102 21158
rect 7603 18737 7797 21903
rect 8234 19006 8445 22535
rect 8882 19298 9078 23162
rect 9496 19704 9704 23896
rect 10127 20093 10313 24893
rect 10127 19907 10693 20093
rect 9496 19496 10304 19704
rect 8882 19102 9638 19298
rect 8234 18795 9045 19006
rect 7603 18543 8437 18737
rect 8243 18497 8437 18543
rect 6898 18238 7658 18442
rect 7862 18238 7868 18442
rect 8243 18297 8437 18303
rect 8834 18506 9045 18795
rect 9442 18498 9638 19102
rect 9442 18296 9638 18302
rect 10096 18504 10304 19496
rect 10507 18493 10693 19907
rect 10507 18307 10707 18493
rect 10893 18307 10899 18493
rect 11339 18477 11493 24877
rect 12547 22465 12677 24865
rect 11935 22335 12677 22465
rect 11935 18465 12065 22335
rect 13700 21938 13916 24808
rect 11935 18329 12065 18335
rect 12572 21722 13916 21938
rect 12572 18498 12788 21722
rect 11339 18317 11493 18323
rect 8834 18289 9045 18295
rect 10096 18290 10304 18296
rect 12572 18276 12788 18282
rect 14024 20785 14216 20786
rect 14910 20785 15099 24675
rect 14024 20596 15099 20785
rect 16099 20782 16302 24772
rect 17299 21947 17493 24807
rect 23631 21947 23829 21949
rect 17299 21753 23829 21947
rect 14024 18466 14216 20596
rect 16099 20579 21831 20782
rect 21628 18492 21831 20579
rect 23631 19159 23829 21753
rect 23631 18955 23829 18961
rect 14760 18375 15160 18380
rect 14024 18268 14216 18274
rect 14756 17985 14765 18375
rect 15155 17985 15164 18375
rect 22420 18395 22820 18400
rect 21628 18283 21831 18289
rect 22416 18005 22425 18395
rect 22815 18005 22824 18395
rect 6100 17884 6660 17890
rect 14760 17840 15160 17985
rect 14760 17434 15160 17440
rect 22420 17840 22820 18005
rect 22420 17434 22820 17440
rect 21100 13220 21540 13260
rect 15860 13180 16300 13190
rect 15840 12900 15860 13180
rect 16300 12900 16360 13180
rect 15840 12860 16360 12900
rect 15840 12680 15860 12860
rect 16300 12680 16360 12860
rect 15840 12660 16360 12680
rect 21100 12960 21160 13220
rect 21480 12960 21540 13220
rect 21100 12920 21540 12960
rect 21100 12660 21160 12920
rect 21480 12660 21540 12920
rect 21160 12650 21480 12660
rect 16240 10480 16700 10820
rect 16900 9420 18860 9440
rect 16900 9320 16960 9420
rect 18740 9320 18860 9420
rect 16900 9280 18860 9320
rect 16900 9140 16960 9280
rect 18740 9140 18860 9280
rect 21740 9360 22400 9380
rect 21740 9260 21780 9360
rect 22360 9260 22400 9360
rect 21740 9240 22400 9260
rect 21740 9200 21780 9240
rect 16900 9100 18860 9140
rect 22360 9200 22400 9240
rect 21780 9130 22360 9140
rect 26216 8069 26624 8073
rect 25665 7651 25671 8069
rect 26089 8064 26629 8069
rect 26089 7656 26216 8064
rect 26624 7656 26629 8064
rect 26089 7651 26629 7656
rect 26216 7647 26624 7651
rect 13980 4400 14860 4420
rect 13980 4100 14020 4400
rect 14240 4380 14860 4400
rect 14240 4120 14500 4380
rect 14820 4120 14860 4380
rect 14240 4100 14860 4120
rect 13980 4080 14860 4100
rect 12000 3860 12320 3940
rect 12000 3620 12040 3860
rect 12300 3620 12320 3860
rect 12000 3608 12320 3620
rect 6420 3200 7020 3240
rect 6420 3060 6460 3200
rect 6980 3060 7020 3200
rect 6420 2920 7020 3060
rect 6420 2740 6460 2920
rect 6980 2740 7020 2920
rect 6420 2720 7020 2740
rect 11972 768 12348 3608
rect 9092 720 12348 768
rect 15340 760 15700 4880
rect 17880 4360 18280 4380
rect 17880 4120 17920 4360
rect 18240 4120 18280 4360
rect 22380 4320 22700 4340
rect 22380 4160 22400 4320
rect 22500 4160 22700 4320
rect 24520 4160 24820 4300
rect 22380 4140 22700 4160
rect 15877 2916 16235 2964
rect 15875 2655 15881 2916
rect 16232 2655 16238 2916
rect 15877 2619 16235 2655
rect 15868 2261 15877 2619
rect 16129 2261 16235 2619
rect 9092 440 9140 720
rect 9440 440 12348 720
rect 9092 392 12348 440
rect 13560 720 15700 760
rect 13560 420 13580 720
rect 13900 420 15700 720
rect 13560 400 15700 420
rect 17880 680 18280 4120
rect 24683 3693 24817 4160
rect 21500 3260 21960 3280
rect 21500 3000 21540 3260
rect 21900 3000 21960 3260
rect 21500 2780 21960 3000
rect 24685 2992 24816 3693
rect 25360 3280 25920 3320
rect 25360 3000 25400 3280
rect 25860 3000 25920 3280
rect 24658 2861 24842 2992
rect 21500 2480 21540 2780
rect 21900 2480 21960 2780
rect 21500 2400 21960 2480
rect 22400 2720 24871 2861
rect 22400 2440 22420 2720
rect 22620 2620 24871 2720
rect 25360 2640 25920 3000
rect 22620 2440 22641 2620
rect 22400 2400 22641 2440
rect 25360 2440 25400 2640
rect 25860 2440 25920 2640
rect 25360 2400 25920 2440
rect 17880 440 17920 680
rect 18240 440 18280 680
rect 17880 400 18280 440
rect 26760 940 27100 980
rect 26760 700 26800 940
rect 27060 700 27100 940
rect 26760 680 27100 700
rect 26760 440 26800 680
rect 27060 440 27100 680
rect 26760 400 27100 440
rect 31260 960 31580 980
rect 31260 680 31280 960
rect 31540 680 31580 960
rect 31260 640 31580 680
rect 31260 440 31280 640
rect 31540 440 31580 640
rect 31260 420 31580 440
<< via2 >>
rect 12558 44898 12641 44981
rect 4191 43470 4290 43569
rect 13305 44725 13374 44794
rect 14044 44584 14115 44655
rect 14765 44445 14835 44515
rect 15498 44278 15581 44361
rect 16236 44076 16324 44164
rect 16984 43884 17057 43957
rect 17724 43744 17795 43815
rect 28016 43596 28103 43683
rect 28733 43313 28827 43407
rect 29497 42817 29583 42903
rect 27282 41998 27366 42082
rect 30953 41653 31047 41747
rect 1200 17890 1760 18450
rect 14765 17985 15155 18375
rect 22425 18005 22815 18395
rect 15860 12900 16300 13180
rect 21160 12960 21480 13220
rect 16960 9140 18740 9280
rect 21780 9140 22360 9240
rect 26216 7656 26624 8064
rect 14500 4120 14820 4380
rect 6460 2740 6980 2920
rect 17920 4120 18240 4360
rect 22400 4160 22500 4320
rect 15877 2261 16129 2619
rect 9140 440 9440 720
rect 13580 420 13900 720
rect 21540 2480 21900 2780
rect 22420 2440 22620 2720
rect 25400 2440 25860 2640
rect 17920 440 18240 680
rect 26800 440 27060 680
rect 31280 440 31540 640
<< metal3 >>
rect 12553 44981 12646 44986
rect 12553 44898 12558 44981
rect 12641 44898 12646 44981
rect 16979 44901 17062 44902
rect 12553 44893 12646 44898
rect 13305 44894 13374 44900
rect 760 44812 9060 44860
rect 760 44748 796 44812
rect 860 44748 1532 44812
rect 1596 44748 2268 44812
rect 2332 44748 3004 44812
rect 3068 44748 3740 44812
rect 3804 44748 4476 44812
rect 4540 44748 5212 44812
rect 5276 44748 5948 44812
rect 6012 44748 6684 44812
rect 6748 44748 7420 44812
rect 7484 44748 8156 44812
rect 8220 44748 8892 44812
rect 8956 44748 9060 44812
rect 760 44720 9060 44748
rect 9520 44812 11220 44860
rect 9520 44748 9628 44812
rect 9692 44748 10364 44812
rect 10428 44748 11100 44812
rect 11164 44748 11220 44812
rect 9520 44720 11220 44748
rect 11818 44842 11903 44848
rect 11818 43680 11903 44757
rect 12558 44842 12641 44893
rect 13305 44799 13374 44825
rect 14044 44895 14115 44901
rect 12558 44753 12641 44759
rect 13300 44794 13379 44799
rect 13300 44725 13305 44794
rect 13374 44725 13379 44794
rect 13300 44720 13379 44725
rect 14044 44660 14115 44824
rect 14765 44895 14835 44901
rect 16236 44884 16324 44890
rect 14039 44655 14120 44660
rect 14039 44584 14044 44655
rect 14115 44584 14120 44655
rect 14039 44579 14120 44584
rect 14765 44520 14835 44825
rect 15498 44861 15581 44867
rect 14760 44515 14840 44520
rect 14760 44445 14765 44515
rect 14835 44445 14840 44515
rect 14760 44440 14840 44445
rect 15498 44366 15581 44778
rect 16974 44820 16980 44901
rect 17061 44820 17067 44901
rect 17724 44895 17795 44901
rect 27277 44826 27371 44827
rect 15493 44361 15586 44366
rect 15493 44278 15498 44361
rect 15581 44278 15586 44361
rect 15493 44273 15586 44278
rect 16236 44169 16324 44796
rect 16231 44164 16329 44169
rect 16231 44076 16236 44164
rect 16324 44076 16329 44164
rect 16231 44071 16329 44076
rect 16979 43957 17062 44820
rect 16979 43884 16984 43957
rect 17057 43884 17062 43957
rect 16979 43879 17062 43884
rect 17724 43820 17795 44824
rect 27272 44734 27278 44826
rect 27370 44734 27376 44826
rect 28016 44803 28103 44809
rect 17719 43815 17800 43820
rect 17719 43744 17724 43815
rect 17795 43744 17800 43815
rect 17719 43739 17800 43744
rect 11818 43580 11900 43680
rect 4180 43569 11900 43580
rect 4180 43470 4191 43569
rect 4290 43470 11900 43569
rect 4180 43460 11900 43470
rect 9617 42623 9704 42624
rect 9612 42538 9618 42623
rect 9703 42538 9709 42623
rect 5320 42140 5640 42180
rect 5310 41900 5320 42140
rect 5640 41900 5650 42140
rect 5320 39440 5640 41900
rect 9617 39864 9704 42538
rect 11320 42140 11640 42180
rect 11310 41900 11320 42140
rect 11640 41900 11650 42140
rect 27277 42082 27371 44734
rect 28016 43688 28103 44716
rect 28733 44807 28827 44813
rect 28011 43683 28108 43688
rect 28011 43596 28016 43683
rect 28103 43596 28108 43683
rect 28011 43591 28108 43596
rect 28733 43412 28827 44713
rect 29497 44803 29583 44809
rect 28728 43407 28832 43412
rect 28728 43313 28733 43407
rect 28827 43313 28832 43407
rect 28728 43308 28832 43313
rect 29497 42908 29583 44717
rect 30953 44767 31047 44827
rect 29492 42903 29588 42908
rect 29492 42817 29497 42903
rect 29583 42817 29588 42903
rect 29492 42812 29588 42817
rect 27277 41998 27282 42082
rect 27366 41998 27371 42082
rect 27277 41993 27371 41998
rect 9617 39771 9704 39777
rect 5320 39280 5360 39440
rect 5600 39280 5640 39440
rect 5320 39260 5640 39280
rect 11320 39440 11640 41900
rect 30953 41752 31047 44673
rect 30948 41747 31052 41752
rect 30948 41653 30953 41747
rect 31047 41653 31052 41747
rect 30948 41648 31052 41653
rect 11320 39280 11360 39440
rect 11600 39280 11640 39440
rect 20451 39397 20457 39483
rect 20543 39397 21677 39483
rect 21763 39397 23777 39483
rect 23863 39397 25377 39483
rect 25463 39397 25523 39483
rect 11320 39260 11640 39280
rect 25397 38363 25483 39397
rect 25397 38271 25483 38277
rect 24217 34886 24344 34887
rect 24075 34761 24081 34886
rect 24479 34761 24485 34886
rect 24217 33304 24344 34761
rect 24217 33171 24344 33177
rect 25355 30245 25485 30251
rect 25355 28545 25485 30115
rect 25355 28409 25485 28415
rect 5300 26560 5640 26596
rect 5300 26360 5320 26560
rect 5620 26360 5640 26560
rect 5300 23360 5640 26360
rect 5300 23040 5320 23360
rect 5620 23040 5640 23360
rect 5300 23020 5640 23040
rect 11300 26580 11640 26620
rect 11300 26380 11320 26580
rect 11620 26380 11640 26580
rect 11300 23360 11640 26380
rect 25775 25346 25904 25351
rect 25774 25345 31074 25346
rect 25774 25216 25775 25345
rect 25904 25216 31074 25345
rect 25774 25215 31074 25216
rect 31205 25215 31211 25346
rect 25775 25210 25904 25215
rect 11300 23040 11320 23360
rect 11620 23040 11640 23360
rect 11300 23020 11640 23040
rect 14760 19839 15160 19840
rect 22420 19839 22820 19840
rect 14755 19441 14761 19839
rect 15159 19441 15165 19839
rect 22415 19441 22421 19839
rect 22819 19441 22825 19839
rect 1195 18450 1765 18455
rect 354 17890 360 18450
rect 920 17890 1200 18450
rect 1760 17890 1765 18450
rect 14760 18375 15160 19441
rect 14760 17985 14765 18375
rect 15155 17985 15160 18375
rect 22420 18395 22820 19441
rect 22420 18005 22425 18395
rect 22815 18005 22820 18395
rect 22420 18000 22820 18005
rect 14760 17980 15160 17985
rect 1195 17885 1765 17890
rect 15840 13540 16360 13600
rect 15840 13260 15880 13540
rect 16320 13260 16360 13540
rect 15840 13180 16360 13260
rect 15840 12900 15860 13180
rect 16300 12900 16360 13180
rect 21100 13540 21540 13600
rect 21100 13280 21160 13540
rect 21480 13280 21540 13540
rect 21100 13220 21540 13280
rect 21100 12960 21160 13220
rect 21480 12960 21540 13220
rect 21100 12920 21540 12960
rect 15840 12860 16360 12900
rect 16260 10660 16680 10920
rect 16840 9280 18860 9320
rect 16840 9140 16960 9280
rect 18740 9140 18860 9280
rect 16840 9100 18860 9140
rect 16840 8960 16960 9100
rect 18740 8960 18860 9100
rect 16840 8880 18860 8960
rect 21740 9240 22380 9300
rect 21740 9140 21780 9240
rect 22360 9140 22380 9240
rect 21740 9060 22380 9140
rect 21740 8960 21780 9060
rect 22360 8960 22380 9060
rect 21740 8940 22380 8960
rect 26892 8069 27308 8074
rect 26211 8068 27309 8069
rect 26211 8064 26892 8068
rect 26211 7656 26216 8064
rect 26624 7656 26892 8064
rect 26211 7652 26892 7656
rect 27308 7652 27309 8068
rect 26211 7651 27309 7652
rect 26892 7646 27308 7651
rect 14479 4380 21411 4411
rect 14479 4120 14500 4380
rect 14820 4360 21411 4380
rect 14820 4120 17920 4360
rect 18240 4340 21411 4360
rect 18240 4320 22520 4340
rect 18240 4160 22400 4320
rect 22500 4160 22520 4320
rect 18240 4120 21411 4160
rect 22390 4155 22510 4160
rect 14479 4089 21411 4120
rect 6420 2920 7020 2960
rect 6420 2740 6460 2920
rect 6980 2740 7020 2920
rect 6420 2340 7020 2740
rect 21500 2780 21960 2880
rect 6420 2060 6460 2340
rect 6980 2060 7020 2340
rect 6420 2020 7020 2060
rect 15808 2619 16198 2635
rect 15808 2261 15877 2619
rect 16129 2395 16198 2619
rect 21500 2480 21540 2780
rect 21900 2480 21960 2780
rect 16129 2261 16395 2395
rect 15808 2005 16395 2261
rect 21500 2340 21960 2480
rect 21500 2060 21540 2340
rect 21900 2060 21960 2340
rect 21500 2020 21960 2060
rect 22340 2720 22680 2780
rect 22340 2440 22420 2720
rect 22620 2440 22680 2720
rect 9100 720 9460 760
rect 9100 440 9140 720
rect 9440 440 9460 720
rect 9100 380 9460 440
rect 9100 180 9140 380
rect 9420 180 9460 380
rect 9100 140 9460 180
rect 13560 720 13920 760
rect 13560 420 13580 720
rect 13900 420 13920 720
rect 13560 380 13920 420
rect 13560 180 13580 380
rect 13900 180 13920 380
rect 13560 160 13920 180
rect 17880 680 18280 700
rect 17880 440 17920 680
rect 18240 440 18280 680
rect 17880 420 18280 440
rect 17880 180 17920 420
rect 18240 180 18280 420
rect 22340 440 22680 2440
rect 25360 2640 25920 2660
rect 25360 2440 25400 2640
rect 25860 2440 25920 2640
rect 25360 2320 25920 2440
rect 25360 2080 25400 2320
rect 25860 2080 25920 2320
rect 25360 2040 25920 2080
rect 22340 260 22420 440
rect 22620 260 22680 440
rect 26760 680 27100 700
rect 26760 440 26800 680
rect 27060 440 27100 680
rect 26760 380 27100 440
rect 22400 220 22640 260
rect 26760 240 26800 380
rect 27040 240 27100 380
rect 26760 200 27100 240
rect 31260 640 31580 660
rect 31260 440 31280 640
rect 31540 440 31580 640
rect 31260 400 31580 440
rect 31260 240 31280 400
rect 31540 240 31580 400
rect 31260 220 31580 240
rect 17880 120 18280 180
<< via3 >>
rect 796 44748 860 44812
rect 1532 44748 1596 44812
rect 2268 44748 2332 44812
rect 3004 44748 3068 44812
rect 3740 44748 3804 44812
rect 4476 44748 4540 44812
rect 5212 44748 5276 44812
rect 5948 44748 6012 44812
rect 6684 44748 6748 44812
rect 7420 44748 7484 44812
rect 8156 44748 8220 44812
rect 8892 44748 8956 44812
rect 9628 44748 9692 44812
rect 10364 44748 10428 44812
rect 11100 44748 11164 44812
rect 11818 44757 11903 44842
rect 12558 44759 12641 44842
rect 13305 44825 13374 44894
rect 14044 44824 14115 44895
rect 14765 44825 14835 44895
rect 15498 44778 15581 44861
rect 16236 44796 16324 44884
rect 16980 44820 17061 44901
rect 17724 44824 17795 44895
rect 27278 44734 27370 44826
rect 9618 42538 9703 42623
rect 5320 41900 5640 42140
rect 11320 41900 11640 42140
rect 28016 44716 28103 44803
rect 28733 44713 28827 44807
rect 29497 44717 29583 44803
rect 30953 44673 31047 44767
rect 9617 39777 9704 39864
rect 5360 39280 5600 39440
rect 11360 39280 11600 39440
rect 20457 39397 20543 39483
rect 21677 39397 21763 39483
rect 23777 39397 23863 39483
rect 25377 39397 25463 39483
rect 25397 38277 25483 38363
rect 24081 34761 24479 34886
rect 24217 33177 24344 33304
rect 25355 30115 25485 30245
rect 25355 28415 25485 28545
rect 5320 26360 5620 26560
rect 5320 23040 5620 23360
rect 11320 26380 11620 26580
rect 25775 25216 25904 25345
rect 31074 25215 31205 25346
rect 11320 23040 11620 23360
rect 14761 19441 15159 19839
rect 22421 19441 22819 19839
rect 360 17890 920 18450
rect 15880 13260 16320 13540
rect 21160 13280 21480 13540
rect 16960 8960 18740 9100
rect 21780 8960 22360 9060
rect 26892 7652 27308 8068
rect 6460 2060 6980 2340
rect 21540 2060 21900 2340
rect 9140 180 9420 380
rect 13580 180 13900 380
rect 17920 180 18240 420
rect 25400 2080 25860 2320
rect 22420 260 22620 440
rect 26800 240 27040 380
rect 31280 240 31540 400
<< metal4 >>
rect 798 44813 858 45152
rect 1534 44813 1594 45152
rect 2270 44813 2330 45152
rect 3006 44813 3066 45152
rect 3742 44813 3802 45152
rect 4478 44813 4538 45152
rect 5214 44813 5274 45152
rect 5950 44813 6010 45152
rect 6686 44813 6746 45152
rect 7422 44813 7482 45152
rect 8158 45150 8218 45152
rect 795 44812 861 44813
rect 795 44748 796 44812
rect 860 44748 861 44812
rect 795 44747 861 44748
rect 1531 44812 1597 44813
rect 1531 44748 1532 44812
rect 1596 44748 1597 44812
rect 1531 44747 1597 44748
rect 2267 44812 2333 44813
rect 2267 44748 2268 44812
rect 2332 44748 2333 44812
rect 2267 44747 2333 44748
rect 3003 44812 3069 44813
rect 3003 44748 3004 44812
rect 3068 44748 3069 44812
rect 3003 44747 3069 44748
rect 3739 44812 3805 44813
rect 3739 44748 3740 44812
rect 3804 44748 3805 44812
rect 3739 44747 3805 44748
rect 4475 44812 4541 44813
rect 4475 44748 4476 44812
rect 4540 44748 4541 44812
rect 4475 44747 4541 44748
rect 5211 44812 5277 44813
rect 5211 44748 5212 44812
rect 5276 44748 5277 44812
rect 5211 44747 5277 44748
rect 5947 44812 6013 44813
rect 5947 44748 5948 44812
rect 6012 44748 6013 44812
rect 5947 44747 6013 44748
rect 6683 44812 6749 44813
rect 6683 44748 6684 44812
rect 6748 44748 6749 44812
rect 6683 44747 6749 44748
rect 7419 44812 7485 44813
rect 7419 44748 7420 44812
rect 7484 44748 7485 44812
rect 7419 44747 7485 44748
rect 8140 44812 8260 45150
rect 8894 44813 8954 45152
rect 9630 45150 9690 45152
rect 8140 44748 8156 44812
rect 8220 44748 8260 44812
rect 8140 44720 8260 44748
rect 8891 44812 8957 44813
rect 8891 44748 8892 44812
rect 8956 44748 8957 44812
rect 8891 44747 8957 44748
rect 9610 44812 9730 45150
rect 10366 44813 10426 45152
rect 11102 45150 11162 45152
rect 11838 45150 11898 45152
rect 12574 45150 12634 45152
rect 13310 45150 13370 45152
rect 14046 45150 14106 45152
rect 14782 45150 14842 45152
rect 15518 45150 15578 45152
rect 16254 45150 16314 45152
rect 16990 45150 17050 45152
rect 17726 45150 17786 45152
rect 18462 45150 18522 45152
rect 9610 44748 9628 44812
rect 9692 44748 9730 44812
rect 9610 44720 9730 44748
rect 10363 44812 10429 44813
rect 10363 44748 10364 44812
rect 10428 44748 10429 44812
rect 10363 44747 10429 44748
rect 11080 44812 11200 45150
rect 11080 44748 11100 44812
rect 11164 44748 11200 44812
rect 11080 44720 11200 44748
rect 11800 44842 11920 45150
rect 11800 44757 11818 44842
rect 11903 44757 11920 44842
rect 11800 44720 11920 44757
rect 12550 44842 12670 45150
rect 12550 44759 12558 44842
rect 12641 44759 12670 44842
rect 12550 44720 12670 44759
rect 13280 44894 13400 45150
rect 13280 44825 13305 44894
rect 13374 44825 13400 44894
rect 13280 44720 13400 44825
rect 14020 44895 14140 45150
rect 14020 44824 14044 44895
rect 14115 44824 14140 44895
rect 14020 44720 14140 44824
rect 14740 44895 14860 45150
rect 14740 44825 14765 44895
rect 14835 44825 14860 44895
rect 14740 44720 14860 44825
rect 15480 44861 15600 45150
rect 15480 44778 15498 44861
rect 15581 44778 15600 44861
rect 15480 44720 15600 44778
rect 16220 44884 16340 45150
rect 16220 44796 16236 44884
rect 16324 44796 16340 44884
rect 16220 44720 16340 44796
rect 16960 44901 17080 45150
rect 16960 44820 16980 44901
rect 17061 44820 17080 44901
rect 16960 44720 17080 44820
rect 17710 44895 17830 45150
rect 18430 44910 18550 45150
rect 17710 44824 17724 44895
rect 17795 44824 17830 44895
rect 17710 44720 17830 44824
rect 18429 44809 18550 44910
rect 19198 44820 19258 45152
rect 19934 44820 19994 45152
rect 20670 44820 20730 45152
rect 21406 44820 21466 45152
rect 22142 44820 22202 45152
rect 22878 44820 22938 45152
rect 23614 44820 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 45150 27354 45152
rect 28030 45150 28090 45152
rect 28766 45150 28826 45152
rect 29502 45150 29562 45152
rect 30238 45150 30298 45152
rect 30974 45150 31034 45152
rect 31710 45150 31770 45152
rect 27260 44826 27380 45150
rect 18430 44720 18550 44809
rect 27260 44734 27278 44826
rect 27370 44734 27380 44826
rect 27260 44720 27380 44734
rect 28000 44803 28120 45150
rect 28000 44720 28016 44803
rect 200 39960 500 44552
rect 8140 42260 8237 44720
rect 9617 42623 9704 44720
rect 28015 44716 28016 44720
rect 28103 44720 28120 44803
rect 28730 44807 28850 45150
rect 28730 44720 28733 44807
rect 28103 44716 28104 44720
rect 28015 44715 28104 44716
rect 28732 44713 28733 44720
rect 28827 44720 28850 44807
rect 29480 44803 29600 45150
rect 29480 44720 29497 44803
rect 28827 44713 28828 44720
rect 29496 44717 29497 44720
rect 29583 44720 29600 44803
rect 30220 44720 30340 45150
rect 30950 44767 31050 45150
rect 31690 44940 31790 45150
rect 30950 44730 30953 44767
rect 29583 44717 29584 44720
rect 29496 44716 29584 44717
rect 28732 44712 28828 44713
rect 30952 44673 30953 44730
rect 31047 44730 31050 44767
rect 31047 44673 31048 44730
rect 30952 44672 31048 44673
rect 9617 42538 9618 42623
rect 9703 42538 9704 42623
rect 9617 42537 9704 42538
rect 31000 42260 31300 44552
rect 5260 42140 31320 42260
rect 5260 41900 5320 42140
rect 5640 41900 11320 42140
rect 11640 41900 31320 42140
rect 5260 41860 31320 41900
rect 200 39864 18700 39960
rect 200 39777 9617 39864
rect 9704 39777 18700 39864
rect 200 39560 18700 39777
rect 200 26100 500 39560
rect 2860 26100 3180 39560
rect 5320 39440 5620 39480
rect 5320 39280 5360 39440
rect 5600 39280 5620 39440
rect 5320 37940 5620 39280
rect 6020 37360 6420 39560
rect 11320 39440 11640 39460
rect 11320 39280 11360 39440
rect 11600 39280 11640 39440
rect 11320 37920 11640 39280
rect 12040 37360 12440 39560
rect 5300 26560 5640 28296
rect 5300 26420 5320 26560
rect 5319 26360 5320 26420
rect 5620 26420 5640 26560
rect 5620 26360 5621 26420
rect 5319 26359 5621 26360
rect 6040 26100 6380 26780
rect 11300 26580 11640 28296
rect 11300 26420 11320 26580
rect 11319 26380 11320 26420
rect 11620 26420 11640 26580
rect 11620 26380 11621 26420
rect 11319 26379 11621 26380
rect 12040 26100 12380 27692
rect 18380 26100 18700 39560
rect 200 25700 18700 26100
rect 20320 39483 20640 41860
rect 21660 40900 22540 40940
rect 20320 39397 20457 39483
rect 20543 39397 20640 39483
rect 21620 40740 22600 40900
rect 23400 40880 24340 40920
rect 21620 40360 21820 40740
rect 22400 40360 22600 40740
rect 21620 40200 22600 40360
rect 23360 40720 24340 40880
rect 23360 40260 23560 40720
rect 23360 40220 24300 40260
rect 24880 40240 25080 40920
rect 25820 40240 26020 40920
rect 21620 40160 22560 40200
rect 21620 39483 21820 40160
rect 23360 40100 24340 40220
rect 24880 40100 26020 40240
rect 23400 40060 24340 40100
rect 24920 40060 25980 40100
rect 24140 39620 24340 40060
rect 21620 39420 21677 39483
rect 200 18460 500 25700
rect 20320 23400 20640 39397
rect 21676 39397 21677 39420
rect 21763 39420 21820 39483
rect 23360 39483 24340 39620
rect 23360 39420 23777 39483
rect 21763 39397 21764 39420
rect 21676 39396 21764 39397
rect 23776 39397 23777 39420
rect 23863 39460 24340 39483
rect 25340 39483 25540 40060
rect 23863 39420 24300 39460
rect 25340 39420 25377 39483
rect 23863 39397 23864 39420
rect 23776 39396 23864 39397
rect 25376 39397 25377 39420
rect 25463 39420 25540 39483
rect 25463 39397 25464 39420
rect 25376 39396 25464 39397
rect 24280 38363 26880 38480
rect 24280 38280 25397 38363
rect 24080 38277 25397 38280
rect 25483 38280 26880 38363
rect 25483 38277 27080 38280
rect 24080 38080 27080 38277
rect 24080 36880 24480 38080
rect 26680 36880 27080 38080
rect 24080 36480 27080 36880
rect 24080 34886 24480 36480
rect 24080 34761 24081 34886
rect 24479 34761 24480 34886
rect 24080 34680 24480 34761
rect 26680 34680 27080 36480
rect 24080 33464 26680 33640
rect 24080 33337 24217 33464
rect 24344 33337 26680 33464
rect 24080 33304 26680 33337
rect 24080 33177 24217 33304
rect 24344 33240 26680 33304
rect 24344 33177 24480 33240
rect 24080 30440 24480 33177
rect 26280 32840 27080 33240
rect 26680 30840 27080 32840
rect 26280 30440 27080 30840
rect 24080 30245 26680 30440
rect 24080 30115 25355 30245
rect 25485 30115 26680 30245
rect 24080 30040 26680 30115
rect 24680 28545 26480 28680
rect 24680 28480 25355 28545
rect 24480 28415 25355 28480
rect 25485 28480 26480 28545
rect 25485 28415 26680 28480
rect 24480 28280 26680 28415
rect 24280 28080 24880 28280
rect 24080 27880 24880 28080
rect 26280 27880 26880 28280
rect 24080 25880 24480 27880
rect 24080 25680 24880 25880
rect 24280 25480 24880 25680
rect 26280 25480 26880 25880
rect 24480 25345 26680 25480
rect 24480 25216 25775 25345
rect 25904 25280 26680 25345
rect 31000 25346 31300 41860
rect 25904 25216 26480 25280
rect 24480 25080 26480 25216
rect 31000 25215 31074 25346
rect 31205 25215 31300 25346
rect 31000 23400 31300 25215
rect 3900 23360 31300 23400
rect 3900 23040 5320 23360
rect 5620 23040 11320 23360
rect 11620 23040 31300 23360
rect 3900 23000 31300 23040
rect 31000 20120 31300 23000
rect 14760 19839 31300 20120
rect 14760 19441 14761 19839
rect 15159 19720 22421 19839
rect 15159 19441 15160 19720
rect 14760 19440 15160 19441
rect 22420 19441 22421 19720
rect 22819 19720 31300 19839
rect 22819 19441 22820 19720
rect 22420 19440 22820 19441
rect 200 18450 960 18460
rect 200 17890 360 18450
rect 920 17890 960 18450
rect 200 17880 960 17890
rect 200 13600 500 17880
rect 200 13540 22400 13600
rect 200 13260 15880 13540
rect 16320 13280 21160 13540
rect 21480 13280 22400 13540
rect 16320 13260 22400 13280
rect 200 13200 22400 13260
rect 200 9200 500 13200
rect 200 9100 22400 9200
rect 200 8960 16960 9100
rect 18740 9060 22400 9100
rect 18740 8960 21780 9060
rect 22360 8960 22400 9060
rect 200 8800 22400 8960
rect 210 8600 500 8800
rect 200 2400 500 8600
rect 31000 8069 31300 19720
rect 26891 8068 31300 8069
rect 26891 7652 26892 8068
rect 27308 7652 31300 8068
rect 26891 7651 31300 7652
rect 200 2340 25920 2400
rect 200 2060 6460 2340
rect 6980 2060 21540 2340
rect 21900 2320 25920 2340
rect 21900 2080 25400 2320
rect 25860 2080 25920 2320
rect 21900 2060 25920 2080
rect 200 2000 25920 2060
rect 200 1400 500 2000
rect 31000 1400 31300 7651
rect 22400 440 22640 460
rect 9100 380 9460 440
rect 400 0 520 200
rect 4816 0 4936 200
rect 9100 180 9140 380
rect 9420 180 9460 380
rect 9100 0 9460 180
rect 13560 380 13920 430
rect 13560 180 13580 380
rect 13900 180 13920 380
rect 13560 0 13920 180
rect 17880 420 18280 440
rect 22400 430 22420 440
rect 17880 180 17920 420
rect 18240 180 18280 420
rect 17880 0 18280 180
rect 22340 260 22420 430
rect 22620 430 22640 440
rect 22620 260 22700 430
rect 22340 0 22700 260
rect 26760 380 27120 430
rect 26760 240 26800 380
rect 27040 240 27120 380
rect 26760 0 27120 240
rect 31260 400 31620 430
rect 31260 240 31280 400
rect 31540 240 31620 400
rect 31260 0 31620 240
use p3_opamp  p3_opamp_0
timestamp 1713301548
transform 1 0 17840 0 1 -200
box 3650 3170 8500 8260
use wowa_analog  wowa_analog_0
timestamp 1713251032
transform 1 0 1626 0 1 -22900
box 4762 25894 25772 41430
use wowa_digital  wowa_digital_0
timestamp 1713283579
transform 1 0 3366 0 1 24460
box 842 0 14062 17164
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31000 1400 31300 44552 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel space 200 1400 500 44552 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal4 210 43270 500 43780 1 VGND
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
