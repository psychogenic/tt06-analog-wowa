magic
tech sky130A
magscale 1 2
timestamp 1713381503
<< metal1 >>
rect 23560 19159 29606 19206
rect 23560 18961 23631 19159
rect 23829 18961 29606 19159
rect 23560 18873 29606 18961
rect 6094 17890 6100 18450
rect 6660 17890 7300 18450
rect 7658 18442 7862 18448
rect 7538 18238 7658 18442
rect 8237 18303 8243 18497
rect 8437 18303 8443 18497
rect 8828 18295 8834 18506
rect 9045 18295 9051 18506
rect 9436 18302 9442 18498
rect 9638 18302 9644 18498
rect 9896 18296 10096 18504
rect 10304 18296 10310 18504
rect 10707 18493 10893 18499
rect 10507 18307 10707 18493
rect 11333 18323 11339 18477
rect 11493 18323 11499 18477
rect 11929 18335 11935 18465
rect 12065 18335 12071 18465
rect 10707 18301 10893 18307
rect 12566 18282 12572 18498
rect 12788 18282 12794 18498
rect 7658 18232 7862 18238
rect 12572 17942 12788 18282
rect 14018 18274 14024 18466
rect 14216 18274 14222 18466
rect 21622 18289 21628 18492
rect 21831 18289 21837 18492
rect 14024 17944 14216 18274
rect 21628 17929 21831 18289
rect 23586 18260 23867 18873
rect 14754 17440 14760 17840
rect 15160 17440 15166 17840
rect 22414 17440 22420 17840
rect 22820 17440 22826 17840
rect 14760 16640 15160 17440
rect 22420 17080 22820 17440
rect 15850 12680 15860 12860
rect 16300 12680 16310 12860
rect 21150 12660 21160 12920
rect 21480 12660 21490 12920
rect 16950 9320 16960 9420
rect 18740 9320 18750 9420
rect 21770 9260 21780 9360
rect 22360 9260 22370 9360
rect 25671 8069 26089 8075
rect 25671 7645 26089 7651
rect 25744 6924 27120 7277
rect 14010 4100 14020 4400
rect 14240 4100 14250 4400
rect 15360 4060 15700 4540
rect 12030 3620 12040 3860
rect 12300 3620 12310 3860
rect 6450 3060 6460 3200
rect 6980 3060 6990 3200
rect 15910 3116 16202 3286
rect 15881 2916 16232 3116
rect 21530 3000 21540 3260
rect 21900 3000 21910 3260
rect 25390 3000 25400 3280
rect 25860 3000 25870 3280
rect 15881 2565 16232 2655
rect 26752 940 27105 6924
rect 26752 700 26800 940
rect 27060 700 27105 940
rect 26752 644 27105 700
rect 29273 987 29606 18873
rect 29273 983 31366 987
rect 29273 960 31583 983
rect 29273 680 31280 960
rect 31540 680 31583 960
rect 29273 657 31583 680
rect 29273 654 31366 657
<< via1 >>
rect 23631 18961 23829 19159
rect 6100 17890 6660 18450
rect 7658 18238 7862 18442
rect 8243 18303 8437 18497
rect 8834 18295 9045 18506
rect 9442 18302 9638 18498
rect 10096 18296 10304 18504
rect 10707 18307 10893 18493
rect 11339 18323 11493 18477
rect 11935 18335 12065 18465
rect 12572 18282 12788 18498
rect 14024 18274 14216 18466
rect 21628 18289 21831 18492
rect 14760 17440 15160 17840
rect 22420 17440 22820 17840
rect 15860 12680 16300 12860
rect 21160 12660 21480 12920
rect 16960 9320 18740 9420
rect 21780 9260 22360 9360
rect 25671 7651 26089 8069
rect 14020 4100 14240 4400
rect 12040 3620 12300 3860
rect 6460 3060 6980 3200
rect 21540 3000 21900 3260
rect 25400 3000 25860 3280
rect 15881 2655 16232 2916
rect 26800 700 27060 940
rect 31280 680 31540 960
<< metal2 >>
rect 30951 44715 31050 44720
rect 11810 44620 11910 44629
rect 30946 44625 30955 44715
rect 31045 44625 31054 44715
rect 11810 44500 11910 44520
rect 4100 44400 11910 44500
rect 12550 44610 12650 44619
rect 4100 42200 4200 44400
rect 12550 44300 12650 44510
rect 5300 44290 12650 44300
rect 5200 44200 12650 44290
rect 13290 44610 13390 44619
rect 5200 42200 5300 44200
rect 13290 44100 13390 44510
rect 6200 44000 13390 44100
rect 14030 44610 14130 44619
rect 14741 44510 14750 44610
rect 14850 44510 14859 44610
rect 15490 44590 15590 44599
rect 6290 42210 6390 44000
rect 14030 43900 14130 44510
rect 7400 43800 14140 43900
rect 7400 42210 7500 43800
rect 14750 43700 14850 44510
rect 8500 43600 14860 43700
rect 8500 42210 8600 43600
rect 15490 43500 15590 44490
rect 16230 44590 16330 44599
rect 16961 44490 16970 44590
rect 17070 44490 17079 44590
rect 17730 44570 17830 44579
rect 9590 43400 15600 43500
rect 9590 42230 9690 43400
rect 16230 43300 16330 44490
rect 10700 43200 16340 43300
rect 10710 42210 10810 43200
rect 16970 43100 17070 44490
rect 11800 43000 17080 43100
rect 11810 42210 11910 43000
rect 17730 42900 17830 44470
rect 12900 42800 17840 42900
rect 12910 42230 13010 42800
rect 14010 42600 14110 42609
rect 14010 42210 14110 42500
rect 15120 42600 15220 42609
rect 15120 42210 15220 42500
rect 16220 42600 16320 42609
rect 16220 42210 16320 42500
rect 17330 42600 17430 42609
rect 17330 42220 17430 42500
rect 30951 42210 31050 44625
rect 18441 42111 31050 42210
rect 4128 21022 4333 25382
rect 5423 21587 5617 25387
rect 6695 22315 6906 25375
rect 7992 23068 8188 25358
rect 9266 23764 9474 25364
rect 9266 23556 9704 23764
rect 10627 23763 10813 25383
rect 7992 22872 9078 23068
rect 6695 22104 8445 22315
rect 5423 21393 7797 21587
rect 6898 21022 7102 21030
rect 4128 20818 7102 21022
rect 6100 18450 6660 18456
rect 1191 17890 1200 18450
rect 1760 17890 6100 18450
rect 6898 18442 7102 20818
rect 7603 18737 7797 21393
rect 8234 19006 8445 22104
rect 8882 19298 9078 22872
rect 9496 19704 9704 23556
rect 10507 23577 10813 23763
rect 9496 19496 10304 19704
rect 8882 19102 9638 19298
rect 8234 18795 9045 19006
rect 7603 18543 8437 18737
rect 8243 18497 8437 18543
rect 6898 18238 7658 18442
rect 7862 18238 7868 18442
rect 8243 18297 8437 18303
rect 8834 18506 9045 18795
rect 9442 18498 9638 19102
rect 9442 18296 9638 18302
rect 10096 18504 10304 19496
rect 10507 18493 10693 23577
rect 11873 23047 12027 25347
rect 11339 22893 12027 23047
rect 10507 18307 10707 18493
rect 10893 18307 10899 18493
rect 11339 18477 11493 22893
rect 13126 22304 13333 25383
rect 11880 22097 13333 22304
rect 11880 18465 12088 22097
rect 14412 21558 14628 25388
rect 11880 18430 11935 18465
rect 12065 18430 12088 18465
rect 12572 21342 14628 21558
rect 12572 18498 12788 21342
rect 11935 18329 12065 18335
rect 11339 18317 11493 18323
rect 8834 18289 9045 18295
rect 10096 18290 10304 18296
rect 12572 18276 12788 18282
rect 14024 20785 14216 20786
rect 15705 20785 15894 25374
rect 14024 20596 15894 20785
rect 17008 20782 17213 25402
rect 18283 21947 18477 25397
rect 23631 21947 23829 21949
rect 18283 21753 23829 21947
rect 14024 18466 14216 20596
rect 17008 20579 21831 20782
rect 17008 20578 17213 20579
rect 21628 18492 21831 20579
rect 23631 19159 23829 21753
rect 23631 18955 23829 18961
rect 14760 18375 15160 18380
rect 14024 18268 14216 18274
rect 14756 17985 14765 18375
rect 15155 17985 15164 18375
rect 22420 18395 22820 18400
rect 21628 18283 21831 18289
rect 22416 18005 22425 18395
rect 22815 18005 22824 18395
rect 6100 17884 6660 17890
rect 14760 17840 15160 17985
rect 14760 17434 15160 17440
rect 22420 17840 22820 18005
rect 22420 17434 22820 17440
rect 21100 13220 21540 13260
rect 15860 13180 16300 13190
rect 15840 12900 15860 13180
rect 16300 12900 16360 13180
rect 15840 12860 16360 12900
rect 15840 12680 15860 12860
rect 16300 12680 16360 12860
rect 15840 12660 16360 12680
rect 21100 12960 21160 13220
rect 21480 12960 21540 13220
rect 21100 12920 21540 12960
rect 21100 12660 21160 12920
rect 21480 12660 21540 12920
rect 21160 12650 21480 12660
rect 16240 10480 16700 10820
rect 16900 9420 18860 9440
rect 16900 9320 16960 9420
rect 18740 9320 18860 9420
rect 16900 9280 18860 9320
rect 16900 9140 16960 9280
rect 18740 9140 18860 9280
rect 21740 9360 22400 9380
rect 21740 9260 21780 9360
rect 22360 9260 22400 9360
rect 21740 9240 22400 9260
rect 21740 9200 21780 9240
rect 16900 9100 18860 9140
rect 22360 9200 22400 9240
rect 21780 9130 22360 9140
rect 26216 8069 26624 8073
rect 25665 7651 25671 8069
rect 26089 8064 26629 8069
rect 26089 7656 26216 8064
rect 26624 7656 26629 8064
rect 26089 7651 26629 7656
rect 26216 7647 26624 7651
rect 13980 4400 14860 4420
rect 13980 4100 14020 4400
rect 14240 4380 14860 4400
rect 14240 4120 14500 4380
rect 14820 4120 14860 4380
rect 14240 4100 14860 4120
rect 13980 4080 14860 4100
rect 12000 3860 12320 3940
rect 12000 3620 12040 3860
rect 12300 3620 12320 3860
rect 12000 3608 12320 3620
rect 6420 3200 7020 3240
rect 6420 3060 6460 3200
rect 6980 3060 7020 3200
rect 6420 2920 7020 3060
rect 6420 2740 6460 2920
rect 6980 2740 7020 2920
rect 6420 2720 7020 2740
rect 11972 768 12348 3608
rect 9092 720 12348 768
rect 15340 760 15700 4880
rect 17880 4360 18280 4380
rect 17880 4120 17920 4360
rect 18240 4120 18280 4360
rect 22380 4320 22700 4340
rect 22380 4160 22400 4320
rect 22500 4160 22700 4320
rect 24520 4160 24820 4300
rect 22380 4140 22700 4160
rect 15877 2916 16235 2964
rect 15875 2655 15881 2916
rect 16232 2655 16238 2916
rect 15877 2619 16235 2655
rect 15868 2261 15877 2619
rect 16129 2261 16235 2619
rect 9092 440 9140 720
rect 9440 440 12348 720
rect 9092 392 12348 440
rect 13560 720 15700 760
rect 13560 420 13580 720
rect 13900 420 15700 720
rect 13560 400 15700 420
rect 17880 680 18280 4120
rect 24683 3693 24817 4160
rect 21500 3260 21960 3280
rect 21500 3000 21540 3260
rect 21900 3000 21960 3260
rect 21500 2780 21960 3000
rect 24685 2992 24816 3693
rect 25360 3280 25920 3320
rect 25360 3000 25400 3280
rect 25860 3000 25920 3280
rect 24658 2861 24842 2992
rect 21500 2480 21540 2780
rect 21900 2480 21960 2780
rect 21500 2400 21960 2480
rect 22400 2720 24871 2861
rect 22400 2440 22420 2720
rect 22620 2620 24871 2720
rect 25360 2640 25920 3000
rect 22620 2440 22641 2620
rect 22400 2400 22641 2440
rect 25360 2440 25400 2640
rect 25860 2440 25920 2640
rect 25360 2400 25920 2440
rect 17880 440 17920 680
rect 18240 440 18280 680
rect 17880 400 18280 440
rect 26760 940 27100 980
rect 26760 700 26800 940
rect 27060 700 27100 940
rect 26760 680 27100 700
rect 26760 440 26800 680
rect 27060 440 27100 680
rect 26760 400 27100 440
rect 31260 960 31580 980
rect 31260 680 31280 960
rect 31540 680 31580 960
rect 31260 640 31580 680
rect 31260 440 31280 640
rect 31540 440 31580 640
rect 31260 420 31580 440
<< via2 >>
rect 30955 44625 31045 44715
rect 11810 44520 11910 44620
rect 12550 44510 12650 44610
rect 13290 44510 13390 44610
rect 14030 44510 14130 44610
rect 14750 44510 14850 44610
rect 15490 44490 15590 44590
rect 16230 44490 16330 44590
rect 16970 44490 17070 44590
rect 17730 44470 17830 44570
rect 14010 42500 14110 42600
rect 15120 42500 15220 42600
rect 16220 42500 16320 42600
rect 17330 42500 17430 42600
rect 1200 17890 1760 18450
rect 14765 17985 15155 18375
rect 22425 18005 22815 18395
rect 15860 12900 16300 13180
rect 21160 12960 21480 13220
rect 16960 9140 18740 9280
rect 21780 9140 22360 9240
rect 26216 7656 26624 8064
rect 14500 4120 14820 4380
rect 6460 2740 6980 2920
rect 17920 4120 18240 4360
rect 22400 4160 22500 4320
rect 15877 2261 16129 2619
rect 9140 440 9440 720
rect 13580 420 13900 720
rect 21540 2480 21900 2780
rect 22420 2440 22620 2720
rect 25400 2440 25860 2640
rect 17920 440 18240 680
rect 26800 440 27060 680
rect 31280 440 31540 640
<< metal3 >>
rect 30950 44889 31050 44890
rect 760 44812 9060 44860
rect 760 44748 796 44812
rect 860 44748 1532 44812
rect 1596 44748 2268 44812
rect 2332 44748 3004 44812
rect 3068 44748 3740 44812
rect 3804 44748 4476 44812
rect 4540 44748 5212 44812
rect 5276 44748 5948 44812
rect 6012 44748 6684 44812
rect 6748 44748 7420 44812
rect 7484 44748 8156 44812
rect 8220 44748 8892 44812
rect 8956 44748 9060 44812
rect 760 44720 9060 44748
rect 9520 44812 11220 44860
rect 9520 44748 9628 44812
rect 9692 44748 10364 44812
rect 10428 44748 11100 44812
rect 11164 44748 11220 44812
rect 30945 44791 30951 44889
rect 31049 44791 31055 44889
rect 9520 44720 11220 44748
rect 12550 44750 12650 44756
rect 14030 44750 14130 44756
rect 11795 44621 11801 44739
rect 11919 44621 11925 44739
rect 11805 44620 11915 44621
rect 11805 44520 11810 44620
rect 11910 44520 11915 44620
rect 12550 44615 12650 44650
rect 13270 44739 13420 44750
rect 13270 44621 13281 44739
rect 13399 44621 13420 44739
rect 11805 44515 11915 44520
rect 12545 44610 12655 44615
rect 12545 44510 12550 44610
rect 12650 44510 12655 44610
rect 13270 44610 13420 44621
rect 15490 44750 15590 44756
rect 14030 44615 14130 44650
rect 14750 44730 14850 44736
rect 14750 44615 14850 44630
rect 13270 44510 13290 44610
rect 13390 44510 13420 44610
rect 14025 44610 14135 44615
rect 14025 44510 14030 44610
rect 14130 44510 14135 44610
rect 12545 44505 12655 44510
rect 13285 44505 13395 44510
rect 14025 44505 14135 44510
rect 14745 44610 14855 44615
rect 14745 44510 14750 44610
rect 14850 44510 14855 44610
rect 15490 44595 15590 44650
rect 16230 44730 16330 44736
rect 16230 44595 16330 44630
rect 16970 44730 17070 44736
rect 16970 44595 17070 44630
rect 17730 44730 17830 44736
rect 14745 44505 14855 44510
rect 15485 44590 15595 44595
rect 15485 44490 15490 44590
rect 15590 44490 15595 44590
rect 15485 44485 15595 44490
rect 16225 44590 16335 44595
rect 16225 44490 16230 44590
rect 16330 44490 16335 44590
rect 16225 44485 16335 44490
rect 16965 44590 17075 44595
rect 16965 44490 16970 44590
rect 17070 44490 17075 44590
rect 17730 44575 17830 44630
rect 27270 44619 27370 44730
rect 30950 44715 31050 44791
rect 28000 44649 28100 44680
rect 16965 44485 17075 44490
rect 17725 44570 17835 44575
rect 17725 44470 17730 44570
rect 17830 44470 17835 44570
rect 27255 44501 27261 44619
rect 27379 44501 27385 44619
rect 27995 44531 28001 44649
rect 28119 44531 28125 44649
rect 28740 44640 28840 44660
rect 28730 44639 28850 44640
rect 17725 44465 17835 44470
rect 27270 43520 27370 44501
rect 14010 43420 27370 43520
rect 14010 42605 14110 43420
rect 28000 43190 28100 44531
rect 28725 44521 28731 44639
rect 28849 44521 28855 44639
rect 29490 44609 29590 44630
rect 30950 44625 30955 44715
rect 31045 44625 31050 44715
rect 30950 44620 31050 44625
rect 28730 44360 28850 44521
rect 29475 44491 29481 44609
rect 29599 44491 29605 44609
rect 15120 43090 28100 43190
rect 15120 42605 15220 43090
rect 28740 42890 28840 44360
rect 16220 42790 28840 42890
rect 16220 42605 16320 42790
rect 14005 42600 14115 42605
rect 14005 42500 14010 42600
rect 14110 42500 14115 42600
rect 14005 42495 14115 42500
rect 15115 42600 15225 42605
rect 15115 42500 15120 42600
rect 15220 42500 15225 42600
rect 15115 42495 15225 42500
rect 16215 42600 16325 42605
rect 16215 42500 16220 42600
rect 16320 42500 16325 42600
rect 16215 42495 16325 42500
rect 17325 42600 17435 42605
rect 29490 42600 29590 44491
rect 17325 42500 17330 42600
rect 17430 42500 29590 42600
rect 17325 42495 17435 42500
rect 8280 41199 8780 41230
rect 8280 40801 8331 41199
rect 8729 40801 8780 41199
rect 14331 41150 14729 41199
rect 14331 40840 14380 41150
rect 14700 40840 14729 41150
rect 14331 40801 14729 40840
rect 8280 40750 8780 40801
rect 8350 39710 8710 40750
rect 14349 39699 14712 40801
rect 20451 39397 20457 39483
rect 20543 39397 21677 39483
rect 21763 39397 23777 39483
rect 23863 39397 25377 39483
rect 25463 39397 25523 39483
rect 25397 38363 25483 39397
rect 25397 38271 25483 38277
rect 24217 34886 24344 34887
rect 24075 34761 24081 34886
rect 24479 34761 24485 34886
rect 24217 33304 24344 34761
rect 24217 33171 24344 33177
rect 25355 30245 25485 30251
rect 25355 28545 25485 30115
rect 25355 28409 25485 28415
rect 5350 26550 5750 26564
rect 5350 26300 5370 26550
rect 5720 26300 5750 26550
rect 5350 25540 5750 26300
rect 8350 26070 8740 26700
rect 8350 25780 8380 26070
rect 8720 25780 8740 26070
rect 8350 25750 8740 25780
rect 11330 26550 11750 26564
rect 11330 26300 11350 26550
rect 11720 26300 11750 26550
rect 11330 25540 11750 26300
rect 14360 26060 14750 26700
rect 14360 25770 14380 26060
rect 14720 25770 14750 26060
rect 14360 25750 14750 25770
rect 17330 26550 17750 26564
rect 17330 26300 17360 26550
rect 17730 26300 17750 26550
rect 17330 25540 17750 26300
rect 5356 23394 5744 25540
rect 11335 23436 11746 25540
rect 11335 23019 11746 23025
rect 17337 23414 17744 25540
rect 25775 25346 25904 25351
rect 25774 25345 31074 25346
rect 25774 25216 25775 25345
rect 25904 25216 31074 25345
rect 25774 25215 31074 25216
rect 31205 25215 31211 25346
rect 25775 25210 25904 25215
rect 5356 23000 5744 23006
rect 17337 22997 17744 23007
rect 15824 22405 32416501 22748
rect 14760 19839 15160 19840
rect 22420 19839 22820 19840
rect 14755 19441 14761 19839
rect 15159 19441 15165 19839
rect 22415 19441 22421 19839
rect 22819 19441 22825 19839
rect 1195 18450 1765 18455
rect 354 17890 360 18450
rect 920 17890 1200 18450
rect 1760 17890 1765 18450
rect 14760 18375 15160 19441
rect 14760 17985 14765 18375
rect 15155 17985 15160 18375
rect 22420 18395 22820 19441
rect 22420 18005 22425 18395
rect 22815 18005 22820 18395
rect 22420 18000 22820 18005
rect 14760 17980 15160 17985
rect 1195 17885 1765 17890
rect 15840 13540 16360 13600
rect 15840 13260 15880 13540
rect 16320 13260 16360 13540
rect 15840 13180 16360 13260
rect 15840 12900 15860 13180
rect 16300 12900 16360 13180
rect 21100 13540 21540 13600
rect 21100 13280 21160 13540
rect 21480 13280 21540 13540
rect 21100 13220 21540 13280
rect 21100 12960 21160 13220
rect 21480 12960 21540 13220
rect 21100 12920 21540 12960
rect 15840 12860 16360 12900
rect 16260 10660 16680 10920
rect 16840 9280 18860 9320
rect 16840 9140 16960 9280
rect 18740 9140 18860 9280
rect 16840 9100 18860 9140
rect 16840 8960 16960 9100
rect 18740 8960 18860 9100
rect 16840 8880 18860 8960
rect 21740 9240 22380 9300
rect 21740 9140 21780 9240
rect 22360 9140 22380 9240
rect 21740 9060 22380 9140
rect 21740 8960 21780 9060
rect 22360 8960 22380 9060
rect 21740 8940 22380 8960
rect 26892 8069 27308 8074
rect 26211 8068 27309 8069
rect 26211 8064 26892 8068
rect 26211 7656 26216 8064
rect 26624 7656 26892 8064
rect 26211 7652 26892 7656
rect 27308 7652 27309 8068
rect 26211 7651 27309 7652
rect 26892 7646 27308 7651
rect 14479 4380 21411 4411
rect 14479 4120 14500 4380
rect 14820 4360 21411 4380
rect 14820 4120 17920 4360
rect 18240 4340 21411 4360
rect 18240 4320 22520 4340
rect 18240 4160 22400 4320
rect 22500 4160 22520 4320
rect 18240 4120 21411 4160
rect 22390 4155 22510 4160
rect 14479 4089 21411 4120
rect 6420 2920 7020 2960
rect 6420 2740 6460 2920
rect 6980 2740 7020 2920
rect 6420 2340 7020 2740
rect 21500 2780 21960 2880
rect 6420 2060 6460 2340
rect 6980 2060 7020 2340
rect 6420 2020 7020 2060
rect 15808 2619 16198 2635
rect 15808 2261 15877 2619
rect 16129 2395 16198 2619
rect 21500 2480 21540 2780
rect 21900 2480 21960 2780
rect 16129 2261 16395 2395
rect 15808 2005 16395 2261
rect 21500 2340 21960 2480
rect 21500 2060 21540 2340
rect 21900 2060 21960 2340
rect 21500 2020 21960 2060
rect 22340 2720 22680 2780
rect 22340 2440 22420 2720
rect 22620 2440 22680 2720
rect 9100 720 9460 760
rect 9100 440 9140 720
rect 9440 440 9460 720
rect 9100 380 9460 440
rect 9100 180 9140 380
rect 9420 180 9460 380
rect 9100 140 9460 180
rect 13560 720 13920 760
rect 13560 420 13580 720
rect 13900 420 13920 720
rect 13560 380 13920 420
rect 13560 180 13580 380
rect 13900 180 13920 380
rect 13560 160 13920 180
rect 17880 680 18280 700
rect 17880 440 17920 680
rect 18240 440 18280 680
rect 17880 420 18280 440
rect 17880 180 17920 420
rect 18240 180 18280 420
rect 22340 440 22680 2440
rect 25360 2640 25920 2660
rect 25360 2440 25400 2640
rect 25860 2440 25920 2640
rect 25360 2320 25920 2440
rect 25360 2080 25400 2320
rect 25860 2080 25920 2320
rect 25360 2040 25920 2080
rect 22340 260 22420 440
rect 22620 260 22680 440
rect 26760 680 27100 700
rect 26760 440 26800 680
rect 27060 440 27100 680
rect 26760 380 27100 440
rect 22400 220 22640 260
rect 26760 240 26800 380
rect 27040 240 27100 380
rect 26760 200 27100 240
rect 31260 640 31580 660
rect 31260 440 31280 640
rect 31540 440 31580 640
rect 31260 400 31580 440
rect 31260 240 31280 400
rect 31540 240 31580 400
rect 31260 220 31580 240
rect 17880 120 18280 180
<< via3 >>
rect 796 44748 860 44812
rect 1532 44748 1596 44812
rect 2268 44748 2332 44812
rect 3004 44748 3068 44812
rect 3740 44748 3804 44812
rect 4476 44748 4540 44812
rect 5212 44748 5276 44812
rect 5948 44748 6012 44812
rect 6684 44748 6748 44812
rect 7420 44748 7484 44812
rect 8156 44748 8220 44812
rect 8892 44748 8956 44812
rect 9628 44748 9692 44812
rect 10364 44748 10428 44812
rect 11100 44748 11164 44812
rect 30951 44791 31049 44889
rect 11801 44621 11919 44739
rect 12550 44650 12650 44750
rect 13281 44621 13399 44739
rect 14030 44650 14130 44750
rect 14750 44630 14850 44730
rect 15490 44650 15590 44750
rect 16230 44630 16330 44730
rect 16970 44630 17070 44730
rect 17730 44630 17830 44730
rect 27261 44501 27379 44619
rect 28001 44531 28119 44649
rect 28731 44521 28849 44639
rect 29481 44491 29599 44609
rect 8331 40801 8729 41199
rect 14380 40840 14700 41150
rect 20457 39397 20543 39483
rect 21677 39397 21763 39483
rect 23777 39397 23863 39483
rect 25377 39397 25463 39483
rect 25397 38277 25483 38363
rect 24081 34761 24479 34886
rect 24217 33177 24344 33304
rect 25355 30115 25485 30245
rect 25355 28415 25485 28545
rect 5370 26300 5720 26550
rect 8380 25780 8720 26070
rect 11350 26300 11720 26550
rect 14380 25770 14720 26060
rect 17360 26300 17730 26550
rect 5356 23006 5744 23394
rect 11335 23025 11746 23436
rect 25775 25216 25904 25345
rect 31074 25215 31205 25346
rect 17337 23007 17744 23414
rect 14761 19441 15159 19839
rect 22421 19441 22819 19839
rect 360 17890 920 18450
rect 15880 13260 16320 13540
rect 21160 13280 21480 13540
rect 16960 8960 18740 9100
rect 21780 8960 22360 9060
rect 26892 7652 27308 8068
rect 6460 2060 6980 2340
rect 21540 2060 21900 2340
rect 9140 180 9420 380
rect 13580 180 13900 380
rect 17920 180 18240 420
rect 25400 2080 25860 2320
rect 22420 260 22620 440
rect 26800 240 27040 380
rect 31280 240 31540 400
<< metal4 >>
rect 798 44813 858 45152
rect 1534 44813 1594 45152
rect 2270 44813 2330 45152
rect 3006 44813 3066 45152
rect 3742 44813 3802 45152
rect 4478 44813 4538 45152
rect 5214 44813 5274 45152
rect 5950 44813 6010 45152
rect 6686 44813 6746 45152
rect 7422 44813 7482 45152
rect 8158 45150 8218 45152
rect 795 44812 861 44813
rect 795 44748 796 44812
rect 860 44748 861 44812
rect 795 44747 861 44748
rect 1531 44812 1597 44813
rect 1531 44748 1532 44812
rect 1596 44748 1597 44812
rect 1531 44747 1597 44748
rect 2267 44812 2333 44813
rect 2267 44748 2268 44812
rect 2332 44748 2333 44812
rect 2267 44747 2333 44748
rect 3003 44812 3069 44813
rect 3003 44748 3004 44812
rect 3068 44748 3069 44812
rect 3003 44747 3069 44748
rect 3739 44812 3805 44813
rect 3739 44748 3740 44812
rect 3804 44748 3805 44812
rect 3739 44747 3805 44748
rect 4475 44812 4541 44813
rect 4475 44748 4476 44812
rect 4540 44748 4541 44812
rect 4475 44747 4541 44748
rect 5211 44812 5277 44813
rect 5211 44748 5212 44812
rect 5276 44748 5277 44812
rect 5211 44747 5277 44748
rect 5947 44812 6013 44813
rect 5947 44748 5948 44812
rect 6012 44748 6013 44812
rect 5947 44747 6013 44748
rect 6683 44812 6749 44813
rect 6683 44748 6684 44812
rect 6748 44748 6749 44812
rect 6683 44747 6749 44748
rect 7419 44812 7485 44813
rect 7419 44748 7420 44812
rect 7484 44748 7485 44812
rect 7419 44747 7485 44748
rect 8140 44812 8260 45150
rect 8894 44813 8954 45152
rect 9630 45150 9690 45152
rect 8140 44748 8156 44812
rect 8220 44748 8260 44812
rect 8140 44720 8260 44748
rect 8891 44812 8957 44813
rect 8891 44748 8892 44812
rect 8956 44748 8957 44812
rect 8891 44747 8957 44748
rect 9610 44812 9730 45150
rect 10366 44813 10426 45152
rect 11102 45150 11162 45152
rect 11838 45150 11898 45152
rect 12574 45150 12634 45152
rect 13310 45150 13370 45152
rect 14046 45150 14106 45152
rect 14782 45150 14842 45152
rect 15518 45150 15578 45152
rect 16254 45150 16314 45152
rect 16990 45150 17050 45152
rect 17726 45150 17786 45152
rect 18462 45150 18522 45152
rect 9610 44748 9628 44812
rect 9692 44748 9730 44812
rect 9610 44720 9730 44748
rect 10363 44812 10429 44813
rect 10363 44748 10364 44812
rect 10428 44748 10429 44812
rect 10363 44747 10429 44748
rect 11080 44812 11200 45150
rect 11080 44748 11100 44812
rect 11164 44748 11200 44812
rect 11080 44720 11200 44748
rect 11800 44739 11920 45150
rect 12550 44751 12670 45150
rect 200 41200 500 44552
rect 8140 42260 8237 44720
rect 9617 42537 9704 44720
rect 11800 44621 11801 44739
rect 11919 44621 11920 44739
rect 12549 44750 12670 44751
rect 12549 44650 12550 44750
rect 12650 44650 12670 44750
rect 12549 44649 12670 44650
rect 12550 44640 12670 44649
rect 13280 44739 13400 45150
rect 11800 44620 11920 44621
rect 13280 44621 13281 44739
rect 13399 44621 13400 44739
rect 13280 44620 13400 44621
rect 14020 44750 14140 45150
rect 14020 44650 14030 44750
rect 14130 44650 14140 44750
rect 14020 44620 14140 44650
rect 14740 44730 14860 45150
rect 14740 44630 14750 44730
rect 14850 44630 14860 44730
rect 15480 44750 15600 45150
rect 15480 44650 15490 44750
rect 15590 44650 15600 44750
rect 15480 44640 15600 44650
rect 16220 44730 16340 45150
rect 14740 44600 14860 44630
rect 16220 44630 16230 44730
rect 16330 44630 16340 44730
rect 16220 44620 16340 44630
rect 16960 44730 17080 45150
rect 16960 44630 16970 44730
rect 17070 44630 17080 44730
rect 16960 44620 17080 44630
rect 17710 44731 17830 45150
rect 18430 44910 18550 45150
rect 18429 44809 18550 44910
rect 19198 44820 19258 45152
rect 19934 44820 19994 45152
rect 20670 44820 20730 45152
rect 21406 44820 21466 45152
rect 22142 44820 22202 45152
rect 22878 44820 22938 45152
rect 23614 44820 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 45150 27354 45152
rect 28030 45150 28090 45152
rect 28766 45150 28826 45152
rect 29502 45150 29562 45152
rect 30238 45150 30298 45152
rect 30974 45150 31034 45152
rect 31710 45150 31770 45152
rect 18430 44790 18550 44809
rect 17710 44730 17831 44731
rect 17710 44630 17730 44730
rect 17830 44630 17831 44730
rect 17710 44629 17831 44630
rect 17710 44600 17830 44629
rect 27260 44619 27380 45150
rect 27260 44501 27261 44619
rect 27379 44501 27380 44619
rect 28000 44649 28120 45150
rect 28000 44531 28001 44649
rect 28119 44531 28120 44649
rect 28000 44530 28120 44531
rect 28730 44639 28850 45150
rect 28730 44521 28731 44639
rect 28849 44521 28850 44639
rect 28730 44520 28850 44521
rect 29480 44609 29600 45150
rect 30220 44790 30340 45150
rect 30950 44889 31050 45150
rect 31690 44940 31790 45150
rect 30950 44791 30951 44889
rect 31049 44791 31050 44889
rect 30950 44790 31050 44791
rect 27260 44500 27380 44501
rect 29480 44491 29481 44609
rect 29599 44491 29600 44609
rect 29480 44490 29600 44491
rect 31000 42260 31300 44552
rect 5160 41860 31300 42260
rect 8280 41200 8780 41230
rect 200 41199 18700 41200
rect 200 40801 8331 41199
rect 8729 41150 18700 41199
rect 8729 40840 14380 41150
rect 14700 40840 18700 41150
rect 8729 40801 18700 40840
rect 200 40800 18700 40801
rect 200 26100 500 40800
rect 2860 26100 3180 40800
rect 8280 40750 8780 40800
rect 8330 38530 8730 40750
rect 14350 38530 14750 40800
rect 5350 26550 5750 27304
rect 5350 26300 5370 26550
rect 5720 26300 5750 26550
rect 5350 26280 5750 26300
rect 8360 26100 8730 26890
rect 11330 26550 11750 27304
rect 11330 26300 11350 26550
rect 11720 26300 11750 26550
rect 11330 26280 11750 26300
rect 14360 26100 14730 26880
rect 17330 26550 17750 27304
rect 17330 26300 17360 26550
rect 17730 26300 17750 26550
rect 17330 26280 17750 26300
rect 18380 26100 18700 39560
rect 200 26070 18700 26100
rect 200 25780 8380 26070
rect 8720 26060 18700 26070
rect 8720 25780 14380 26060
rect 200 25770 14380 25780
rect 14720 25770 18700 26060
rect 200 25700 18700 25770
rect 20320 39483 20640 41860
rect 21660 40900 22540 40940
rect 20320 39397 20457 39483
rect 20543 39397 20640 39483
rect 21620 40740 22600 40900
rect 23400 40880 24340 40920
rect 21620 40360 21820 40740
rect 22400 40360 22600 40740
rect 21620 40200 22600 40360
rect 23360 40720 24340 40880
rect 23360 40260 23560 40720
rect 23360 40220 24300 40260
rect 24880 40240 25080 40920
rect 25820 40240 26020 40920
rect 21620 40160 22560 40200
rect 21620 39483 21820 40160
rect 23360 40100 24340 40220
rect 24880 40100 26020 40240
rect 23400 40060 24340 40100
rect 24920 40060 25980 40100
rect 24140 39620 24340 40060
rect 21620 39420 21677 39483
rect 200 18460 500 25700
rect 11334 23436 11747 23437
rect 11334 23400 11335 23436
rect 5330 23394 11335 23400
rect 5330 23006 5356 23394
rect 5744 23025 11335 23394
rect 11746 23400 11747 23436
rect 17336 23414 17745 23415
rect 17336 23400 17337 23414
rect 11746 23025 17337 23400
rect 5744 23007 17337 23025
rect 17744 23400 17745 23414
rect 20320 23400 20640 39397
rect 21676 39397 21677 39420
rect 21763 39420 21820 39483
rect 23360 39483 24340 39620
rect 23360 39420 23777 39483
rect 21763 39397 21764 39420
rect 21676 39396 21764 39397
rect 23776 39397 23777 39420
rect 23863 39460 24340 39483
rect 25340 39483 25540 40060
rect 23863 39420 24300 39460
rect 25340 39420 25377 39483
rect 23863 39397 23864 39420
rect 23776 39396 23864 39397
rect 25376 39397 25377 39420
rect 25463 39420 25540 39483
rect 25463 39397 25464 39420
rect 25376 39396 25464 39397
rect 24280 38363 26880 38480
rect 24280 38280 25397 38363
rect 24080 38277 25397 38280
rect 25483 38280 26880 38363
rect 25483 38277 27080 38280
rect 24080 38080 27080 38277
rect 24080 36880 24480 38080
rect 26680 36880 27080 38080
rect 24080 36480 27080 36880
rect 24080 34886 24480 36480
rect 24080 34761 24081 34886
rect 24479 34761 24480 34886
rect 24080 34680 24480 34761
rect 26680 34680 27080 36480
rect 24080 33464 26680 33640
rect 24080 33337 24217 33464
rect 24344 33337 26680 33464
rect 24080 33304 26680 33337
rect 24080 33177 24217 33304
rect 24344 33240 26680 33304
rect 24344 33177 24480 33240
rect 24080 30440 24480 33177
rect 26280 32840 27080 33240
rect 26680 30840 27080 32840
rect 26280 30440 27080 30840
rect 24080 30245 26680 30440
rect 24080 30115 25355 30245
rect 25485 30115 26680 30245
rect 24080 30040 26680 30115
rect 24680 28545 26480 28680
rect 24680 28480 25355 28545
rect 24480 28415 25355 28480
rect 25485 28480 26480 28545
rect 25485 28415 26680 28480
rect 24480 28280 26680 28415
rect 24280 28080 24880 28280
rect 24080 27880 24880 28080
rect 26280 27880 26880 28280
rect 24080 25880 24480 27880
rect 24080 25680 24880 25880
rect 24280 25480 24880 25680
rect 26280 25480 26880 25880
rect 24480 25345 26680 25480
rect 24480 25216 25775 25345
rect 25904 25280 26680 25345
rect 31000 25346 31300 41860
rect 25904 25216 26480 25280
rect 24480 25080 26480 25216
rect 31000 25215 31074 25346
rect 31205 25215 31300 25346
rect 31000 23400 31300 25215
rect 17744 23007 31300 23400
rect 5744 23006 31300 23007
rect 5330 23000 31300 23006
rect 31000 20120 31300 23000
rect 14760 19839 31300 20120
rect 14760 19441 14761 19839
rect 15159 19720 22421 19839
rect 15159 19441 15160 19720
rect 14760 19440 15160 19441
rect 22420 19441 22421 19720
rect 22819 19720 31300 19839
rect 22819 19441 22820 19720
rect 22420 19440 22820 19441
rect 200 18450 960 18460
rect 200 17890 360 18450
rect 920 17890 960 18450
rect 200 17880 960 17890
rect 200 13600 500 17880
rect 200 13540 22400 13600
rect 200 13260 15880 13540
rect 16320 13280 21160 13540
rect 21480 13280 22400 13540
rect 16320 13260 22400 13280
rect 200 13200 22400 13260
rect 200 9200 500 13200
rect 200 9100 22400 9200
rect 200 8960 16960 9100
rect 18740 9060 22400 9100
rect 18740 8960 21780 9060
rect 22360 8960 22400 9060
rect 200 8800 22400 8960
rect 210 8600 500 8800
rect 200 2400 500 8600
rect 31000 8069 31300 19720
rect 26891 8068 31300 8069
rect 26891 7652 26892 8068
rect 27308 7652 31300 8068
rect 26891 7651 31300 7652
rect 200 2340 25920 2400
rect 200 2060 6460 2340
rect 6980 2060 21540 2340
rect 21900 2320 25920 2340
rect 21900 2080 25400 2320
rect 25860 2080 25920 2320
rect 21900 2060 25920 2080
rect 200 2000 25920 2060
rect 200 1400 500 2000
rect 31000 1400 31300 7651
rect 22400 440 22640 460
rect 9100 380 9460 440
rect 400 0 520 200
rect 4816 0 4936 200
rect 9100 180 9140 380
rect 9420 180 9460 380
rect 9100 0 9460 180
rect 13560 380 13920 430
rect 13560 180 13580 380
rect 13900 180 13920 380
rect 13560 0 13920 180
rect 17880 420 18280 440
rect 22400 430 22420 440
rect 17880 180 17920 420
rect 18240 180 18280 420
rect 17880 0 18280 180
rect 22340 260 22420 430
rect 22620 430 22640 440
rect 22620 260 22700 430
rect 22340 0 22700 260
rect 26760 380 27120 430
rect 26760 240 26800 380
rect 27040 240 27120 380
rect 26760 0 27120 240
rect 31260 400 31620 430
rect 31260 240 31280 400
rect 31540 240 31620 400
rect 31260 0 31620 240
use p3_opamp  p3_opamp_0
timestamp 1713301548
transform 1 0 17840 0 1 -200
box 3650 3170 8500 8260
use wowa_analog  wowa_analog_0
timestamp 1713251032
transform 1 0 1626 0 1 -22900
box 4762 25894 25772 41430
use wowa_digital  wowa_digital_0
timestamp 1713335925
transform 1 0 3442 0 1 24500
box 658 0 15075 17864
<< labels >>
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 31000 1400 31300 44552 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
rlabel metal4 210 43270 500 43780 1 VGND
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
rlabel metal4 230 2040 500 2370 1 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
