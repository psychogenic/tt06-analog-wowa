magic
tech sky130A
magscale 1 2
timestamp 1713335925
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 721 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
<< ndiff >>
rect 27 119 79 177
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 47 163 127
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 161 331 177
rect 277 127 287 161
rect 321 127 331 161
rect 277 47 331 127
rect 361 93 413 177
rect 361 59 371 93
rect 405 59 413 93
rect 361 47 413 59
rect 467 93 519 177
rect 467 59 475 93
rect 509 59 519 93
rect 467 47 519 59
rect 549 161 603 177
rect 549 127 559 161
rect 593 127 603 161
rect 549 47 603 127
rect 633 161 695 177
rect 633 127 649 161
rect 683 127 695 161
rect 633 93 695 127
rect 633 59 649 93
rect 683 59 695 93
rect 633 47 695 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
rect 467 485 519 497
rect 467 451 475 485
rect 509 451 519 485
rect 467 417 519 451
rect 467 383 475 417
rect 509 383 519 417
rect 467 297 519 383
rect 549 485 603 497
rect 549 451 559 485
rect 593 451 603 485
rect 549 417 603 451
rect 549 383 559 417
rect 593 383 603 417
rect 549 349 603 383
rect 549 315 559 349
rect 593 315 603 349
rect 549 297 603 315
rect 633 485 695 497
rect 633 451 649 485
rect 683 451 695 485
rect 633 417 695 451
rect 633 383 649 417
rect 683 383 695 417
rect 633 349 695 383
rect 633 315 649 349
rect 683 315 695 349
rect 633 297 695 315
<< ndiffc >>
rect 35 85 69 119
rect 119 127 153 161
rect 203 59 237 93
rect 287 127 321 161
rect 371 59 405 93
rect 475 59 509 93
rect 559 127 593 161
rect 649 127 683 161
rect 649 59 683 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 475 451 509 485
rect 475 383 509 417
rect 559 451 593 485
rect 559 383 593 417
rect 559 315 593 349
rect 649 451 683 485
rect 649 383 683 417
rect 649 315 683 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 79 265 109 297
rect 163 265 193 297
rect 22 249 193 265
rect 247 261 277 297
rect 331 261 361 297
rect 519 261 549 297
rect 603 263 633 297
rect 603 261 669 263
rect 22 215 32 249
rect 66 215 193 249
rect 22 199 193 215
rect 235 249 397 261
rect 235 215 251 249
rect 285 215 347 249
rect 381 215 397 249
rect 235 203 397 215
rect 519 249 669 261
rect 519 215 535 249
rect 569 215 619 249
rect 653 215 669 249
rect 519 203 669 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 203
rect 331 177 361 203
rect 519 177 549 203
rect 603 202 669 203
rect 603 177 633 202
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
<< polycont >>
rect 32 215 66 249
rect 251 215 285 249
rect 347 215 381 249
rect 535 215 569 249
rect 619 215 653 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 509 527
rect 405 451 475 485
rect 371 417 509 451
rect 405 383 475 417
rect 371 367 509 383
rect 543 485 609 493
rect 543 451 559 485
rect 593 451 609 485
rect 543 417 609 451
rect 543 383 559 417
rect 593 383 609 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 543 349 609 383
rect 543 333 559 349
rect 321 315 559 333
rect 593 315 609 349
rect 103 289 609 315
rect 643 485 719 527
rect 643 451 649 485
rect 683 451 719 485
rect 643 417 719 451
rect 643 383 649 417
rect 683 383 719 417
rect 643 349 719 383
rect 643 315 649 349
rect 683 315 719 349
rect 643 289 719 315
rect 18 249 66 265
rect 18 215 32 249
rect 18 199 66 215
rect 103 161 169 289
rect 214 249 432 255
rect 214 215 251 249
rect 285 215 347 249
rect 381 215 432 249
rect 494 249 719 255
rect 494 215 535 249
rect 569 215 619 249
rect 653 215 719 249
rect 18 119 69 157
rect 103 127 119 161
rect 153 127 169 161
rect 271 161 609 181
rect 271 127 287 161
rect 321 127 559 161
rect 593 127 609 161
rect 643 161 719 177
rect 643 127 649 161
rect 683 127 719 161
rect 18 85 35 119
rect 643 93 719 127
rect 69 85 203 93
rect 18 59 203 85
rect 237 59 371 93
rect 405 59 421 93
rect 459 59 475 93
rect 509 59 525 93
rect 459 17 525 59
rect 643 59 649 93
rect 683 59 719 93
rect 643 17 719 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 A
port 7 nsew
flabel locali s 122 153 156 187 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel locali s 122 289 156 323 0 FreeSans 250 0 0 0 Y
port 8 nsew
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B
port 9 nsew
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 B
port 9 nsew
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 B
port 9 nsew
flabel locali s 677 221 711 255 0 FreeSans 250 0 0 0 C
port 6 nsew
flabel locali s 586 221 620 255 0 FreeSans 250 0 0 0 C
port 6 nsew
flabel locali s 494 221 528 255 0 FreeSans 250 0 0 0 C
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 nand3_2
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 401848
string GDS_FILE wowa_digital_ol.gds
string GDS_START 394622
string path 0.000 2.720 3.680 2.720 
<< end >>
