magic
tech sky130A
magscale 1 2
timestamp 1713137925
<< metal1 >>
rect -40 3710 160 3910
rect 620 3740 3445 3910
rect -550 3570 170 3610
rect -550 3440 -200 3570
rect -50 3440 170 3570
rect 2160 3480 2360 3486
rect -550 3410 170 3440
rect -280 3110 240 3310
rect 1760 3280 2160 3480
rect 2360 3280 2820 3480
rect 2160 3274 2360 3280
rect -550 2750 -350 3030
rect -550 2620 -530 2750
rect -380 2620 -350 2750
rect 1160 2740 1310 3000
rect -550 2590 -350 2620
rect 610 2610 870 2620
rect 1348 2614 1354 2826
rect 1566 2614 1572 2826
rect -278 2248 -272 2432
rect -88 2340 -82 2432
rect 610 2380 620 2610
rect 850 2380 870 2610
rect 2260 2496 2444 2644
rect 2620 2580 2820 3280
rect 2900 3297 3100 3310
rect 2900 3090 3135 3297
rect 2920 2985 3135 3090
rect 2914 2830 2920 2985
rect 3135 2830 3141 2985
rect 2920 2820 3140 2830
rect 3275 2575 3445 3740
rect 610 2360 870 2380
rect 2935 2405 3445 2575
rect -88 2248 140 2340
rect -272 2108 140 2248
rect -260 2100 140 2108
rect -40 1850 160 2050
rect 790 1870 1270 2220
rect 2030 2090 2280 2100
rect 2030 1870 2040 2090
rect 2270 1870 2280 2090
rect 2935 2015 3105 2405
rect 2030 1860 2280 1870
<< via1 >>
rect -200 3440 -50 3570
rect 2160 3280 2360 3480
rect -530 2620 -380 2750
rect 1354 2614 1566 2826
rect -272 2248 -88 2432
rect 620 2380 850 2610
rect 2100 2490 2260 2650
rect 2920 2830 3135 2985
rect 2040 1870 2270 2090
<< metal2 >>
rect -215 3580 250 3590
rect -215 3570 50 3580
rect -215 3440 -200 3570
rect -50 3440 50 3570
rect 210 3440 250 3580
rect -215 3420 250 3440
rect 1150 3405 1159 3607
rect 1361 3405 1370 3607
rect 2154 3280 2160 3480
rect 2360 3280 2366 3480
rect 2160 3131 2360 3140
rect 2920 2990 3135 2991
rect 2900 2985 3150 2990
rect 1354 2961 1566 2966
rect 1350 2940 1359 2961
rect 1340 2826 1359 2940
rect 1561 2826 1570 2961
rect -550 2750 -350 2790
rect -550 2620 -530 2750
rect -380 2620 -350 2750
rect -550 2600 -350 2620
rect -272 2607 -88 2612
rect 610 2610 870 2620
rect -550 2590 -530 2600
rect -540 2480 -530 2590
rect -390 2590 -350 2600
rect -390 2480 -370 2590
rect -540 2470 -370 2480
rect -276 2433 -267 2607
rect -93 2433 -84 2607
rect -272 2432 -88 2433
rect 610 2360 620 2610
rect -272 2242 -88 2248
rect 850 2360 870 2610
rect 1340 2614 1354 2826
rect 1566 2759 1570 2826
rect 2900 2830 2920 2985
rect 3135 2830 3150 2985
rect 2900 2770 3150 2830
rect 1905 2740 2055 2744
rect 1340 2608 1566 2614
rect 1900 2735 2260 2740
rect 1340 2500 1480 2608
rect 1900 2585 1905 2735
rect 2055 2660 2260 2735
rect 2055 2650 2280 2660
rect 2055 2585 2100 2650
rect 1900 2540 2100 2585
rect 2070 2490 2100 2540
rect 2260 2490 2280 2650
rect 2900 2550 2910 2770
rect 3130 2550 3150 2770
rect 2900 2540 3150 2550
rect 2070 2480 2280 2490
rect 620 2236 850 2245
rect 2114 2176 2207 2185
rect 2030 2090 2114 2100
rect 2207 2090 2280 2100
rect 2030 1870 2040 2090
rect 2270 1870 2280 2090
rect 2030 1860 2280 1870
<< via2 >>
rect 50 3440 210 3580
rect 1159 3405 1361 3607
rect 2160 3280 2360 3337
rect 2160 3140 2360 3280
rect 1359 2826 1561 2961
rect -530 2480 -390 2600
rect -267 2433 -93 2607
rect 620 2380 850 2475
rect 620 2245 850 2380
rect 1359 2759 1561 2826
rect 1905 2585 2055 2735
rect 2910 2550 3130 2770
rect 2114 2090 2207 2176
rect 2114 2083 2207 2090
<< metal3 >>
rect 20 3607 1566 3612
rect 20 3580 1159 3607
rect 20 3440 50 3580
rect 210 3440 1159 3580
rect 20 3405 1159 3440
rect 1361 3405 1566 3607
rect 20 3400 1566 3405
rect -272 3011 -88 3012
rect -277 2829 -271 3011
rect -89 2829 -83 3011
rect 1354 2961 1566 3400
rect 2155 3337 2365 3342
rect 2155 3140 2160 3337
rect 2360 3140 2365 3337
rect 2155 3135 2162 3140
rect 2359 3135 2365 3140
rect 2162 2996 2359 3002
rect -540 2750 -370 2770
rect -540 2620 -530 2750
rect -380 2620 -370 2750
rect -540 2600 -370 2620
rect -540 2480 -530 2600
rect -390 2480 -370 2600
rect -540 2470 -370 2480
rect -272 2607 -88 2829
rect 1354 2759 1359 2961
rect 1561 2759 1566 2961
rect 1354 2754 1566 2759
rect 2905 2770 3135 2775
rect 1651 2740 1809 2745
rect -272 2433 -267 2607
rect -93 2433 -88 2607
rect 1650 2739 2060 2740
rect 1650 2581 1651 2739
rect 1809 2735 2060 2739
rect 1809 2585 1905 2735
rect 2055 2585 2060 2735
rect 1809 2581 2060 2585
rect 1650 2580 2060 2581
rect 1651 2575 1809 2580
rect 2905 2550 2910 2770
rect 3130 2550 3135 2770
rect -272 2428 -88 2433
rect 615 2475 855 2480
rect 615 2470 620 2475
rect 850 2470 855 2475
rect 2905 2304 3135 2550
rect 615 2234 855 2240
rect 2114 2246 2207 2252
rect 2109 2083 2114 2181
rect 2207 2083 2212 2181
rect 2109 2078 2212 2083
rect 2900 2076 2906 2304
rect 3134 2076 3140 2304
rect 2905 2075 3135 2076
<< via3 >>
rect -271 2829 -89 3011
rect 2162 3140 2359 3196
rect 2162 3002 2359 3140
rect -530 2620 -380 2750
rect 1651 2581 1809 2739
rect 615 2245 620 2470
rect 620 2245 850 2470
rect 850 2245 855 2470
rect 615 2240 855 2245
rect 2114 2176 2207 2246
rect 2114 2153 2207 2176
rect 2906 2076 3134 2304
<< metal4 >>
rect 2161 3196 2360 3197
rect 2161 3012 2162 3196
rect -272 3011 2162 3012
rect -272 2829 -271 3011
rect -89 3002 2162 3011
rect 2359 3002 2360 3196
rect -89 3001 2360 3002
rect -89 2829 2352 3001
rect -272 2828 2352 2829
rect -540 2750 -290 2770
rect -540 2620 -530 2750
rect -380 2740 -290 2750
rect -380 2739 1810 2740
rect -380 2620 1651 2739
rect -540 2581 1651 2620
rect 1809 2581 1810 2739
rect -540 2580 1810 2581
rect 614 2470 856 2471
rect 614 2240 615 2470
rect 855 2305 856 2470
rect 855 2304 3135 2305
rect 855 2246 2906 2304
rect 855 2240 2114 2246
rect 614 2239 2114 2240
rect 620 2153 2114 2239
rect 2207 2153 2906 2246
rect 620 2076 2906 2153
rect 3134 2076 3135 2304
rect 620 2075 3135 2076
use lvtnot  x1
timestamp 1713131393
transform 1 0 -260 0 1 2580
box 1400 340 2238 1340
use passgate  x2
timestamp 1713131218
transform 0 1 1750 -1 0 4980
box 2200 -700 3200 1400
use passgate  x3
timestamp 1713131218
transform 1 0 -2260 0 1 2510
box 2200 -700 3200 1400
<< labels >>
flabel metal1 2900 3100 3100 3300 0 FreeSans 1280 0 0 0 OUT
port 3 nsew
flabel metal1 -550 2830 -350 3030 0 FreeSans 1280 0 0 0 IN1
port 2 nsew
flabel metal1 -274 3110 -74 3310 0 FreeSans 1280 0 0 0 IN0
port 1 nsew
flabel metal1 -550 3410 -350 3610 0 FreeSans 1280 0 0 0 SEL
port 0 nsew
flabel metal1 -40 3710 160 3910 0 FreeSans 1280 0 0 0 VCC
port 4 nsew
flabel metal1 -40 1850 160 2050 0 FreeSans 1280 0 0 0 VSS
port 5 nsew
rlabel metal1 2360 3280 2820 3480 1 SEL_N
<< end >>
