magic
tech sky130A
magscale 1 2
timestamp 1713335925
<< viali >>
rect 1409 15113 1443 15147
rect 1869 15113 1903 15147
rect 2973 15113 3007 15147
rect 4077 15113 4111 15147
rect 5181 15113 5215 15147
rect 6377 15113 6411 15147
rect 7389 15113 7423 15147
rect 8493 15113 8527 15147
rect 9597 15113 9631 15147
rect 1593 14977 1627 15011
rect 2053 14977 2087 15011
rect 3157 14977 3191 15011
rect 4261 14977 4295 15011
rect 5365 14977 5399 15011
rect 6561 14977 6595 15011
rect 7573 14977 7607 15011
rect 8677 14977 8711 15011
rect 9781 14977 9815 15011
rect 10333 14977 10367 15011
rect 10517 14977 10551 15011
rect 11805 14977 11839 15011
rect 12909 14977 12943 15011
rect 13921 14977 13955 15011
rect 10517 14773 10551 14807
rect 11989 14773 12023 14807
rect 13093 14773 13127 14807
rect 13737 14773 13771 14807
rect 7389 14569 7423 14603
rect 3249 14501 3283 14535
rect 1869 14365 1903 14399
rect 5181 14365 5215 14399
rect 8769 14365 8803 14399
rect 9045 14365 9079 14399
rect 9312 14365 9346 14399
rect 10609 14365 10643 14399
rect 12265 14365 12299 14399
rect 12541 14365 12575 14399
rect 12909 14365 12943 14399
rect 2136 14297 2170 14331
rect 5448 14297 5482 14331
rect 8502 14297 8536 14331
rect 10854 14297 10888 14331
rect 6561 14229 6595 14263
rect 10425 14229 10459 14263
rect 11989 14229 12023 14263
rect 12357 14229 12391 14263
rect 12725 14229 12759 14263
rect 13001 14229 13035 14263
rect 2237 14025 2271 14059
rect 2513 14025 2547 14059
rect 3157 14025 3191 14059
rect 3433 14025 3467 14059
rect 4997 14025 5031 14059
rect 6101 14025 6135 14059
rect 8033 14025 8067 14059
rect 8585 14025 8619 14059
rect 10517 14025 10551 14059
rect 10701 14025 10735 14059
rect 12455 14025 12489 14059
rect 12541 14025 12575 14059
rect 2605 13957 2639 13991
rect 3873 13957 3907 13991
rect 12970 13957 13004 13991
rect 2237 13889 2271 13923
rect 2697 13889 2731 13923
rect 2973 13889 3007 13923
rect 3065 13889 3099 13923
rect 3433 13889 3467 13923
rect 5089 13889 5123 13923
rect 5273 13889 5307 13923
rect 5365 13889 5399 13923
rect 5733 13889 5767 13923
rect 5963 13889 5997 13923
rect 6193 13889 6227 13923
rect 6653 13889 6687 13923
rect 6909 13889 6943 13923
rect 8953 13889 8987 13923
rect 9321 13889 9355 13923
rect 9505 13889 9539 13923
rect 10698 13889 10732 13923
rect 11713 13889 11747 13923
rect 11897 13889 11931 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 12347 13889 12381 13923
rect 12633 13889 12667 13923
rect 3617 13821 3651 13855
rect 8769 13821 8803 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9413 13821 9447 13855
rect 11161 13821 11195 13855
rect 12725 13821 12759 13855
rect 5733 13753 5767 13787
rect 11805 13753 11839 13787
rect 2329 13685 2363 13719
rect 3341 13685 3375 13719
rect 5089 13685 5123 13719
rect 5825 13685 5859 13719
rect 11069 13685 11103 13719
rect 11529 13685 11563 13719
rect 14105 13685 14139 13719
rect 3157 13481 3191 13515
rect 4077 13481 4111 13515
rect 4997 13481 5031 13515
rect 6561 13481 6595 13515
rect 9597 13481 9631 13515
rect 11805 13481 11839 13515
rect 12265 13481 12299 13515
rect 4905 13413 4939 13447
rect 8769 13345 8803 13379
rect 9505 13345 9539 13379
rect 1409 13277 1443 13311
rect 2881 13277 2915 13311
rect 3801 13277 3835 13311
rect 4077 13277 4111 13311
rect 4905 13277 4939 13311
rect 5365 13287 5399 13321
rect 6285 13277 6319 13311
rect 6561 13277 6595 13311
rect 9597 13277 9631 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 1676 13209 1710 13243
rect 3157 13209 3191 13243
rect 8524 13209 8558 13243
rect 2789 13141 2823 13175
rect 2973 13141 3007 13175
rect 3893 13141 3927 13175
rect 5181 13141 5215 13175
rect 5273 13141 5307 13175
rect 6377 13141 6411 13175
rect 7389 13141 7423 13175
rect 9229 13141 9263 13175
rect 1685 12937 1719 12971
rect 5089 12937 5123 12971
rect 6377 12937 6411 12971
rect 9689 12937 9723 12971
rect 11989 12937 12023 12971
rect 12909 12937 12943 12971
rect 13553 12937 13587 12971
rect 4905 12869 4939 12903
rect 6545 12869 6579 12903
rect 6745 12869 6779 12903
rect 9873 12869 9907 12903
rect 1869 12801 1903 12835
rect 8953 12801 8987 12835
rect 9413 12801 9447 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10241 12801 10275 12835
rect 10333 12801 10367 12835
rect 11805 12801 11839 12835
rect 11897 12801 11931 12835
rect 12081 12801 12115 12835
rect 9045 12733 9079 12767
rect 10517 12733 10551 12767
rect 11529 12733 11563 12767
rect 13093 12733 13127 12767
rect 13185 12733 13219 12767
rect 4537 12665 4571 12699
rect 11713 12665 11747 12699
rect 4905 12597 4939 12631
rect 6561 12597 6595 12631
rect 8769 12597 8803 12631
rect 9321 12597 9355 12631
rect 10057 12597 10091 12631
rect 11621 12597 11655 12631
rect 1685 12393 1719 12427
rect 4261 12393 4295 12427
rect 4813 12393 4847 12427
rect 7021 12393 7055 12427
rect 7849 12393 7883 12427
rect 8401 12393 8435 12427
rect 10977 12393 11011 12427
rect 11437 12393 11471 12427
rect 13645 12393 13679 12427
rect 1869 12325 1903 12359
rect 2973 12325 3007 12359
rect 6193 12325 6227 12359
rect 7389 12325 7423 12359
rect 9965 12325 9999 12359
rect 12449 12325 12483 12359
rect 2421 12257 2455 12291
rect 2789 12257 2823 12291
rect 3249 12257 3283 12291
rect 3341 12257 3375 12291
rect 7757 12257 7791 12291
rect 2513 12189 2547 12223
rect 2881 12189 2915 12223
rect 3157 12189 3191 12223
rect 3433 12189 3467 12223
rect 6929 12189 6963 12223
rect 7033 12189 7067 12223
rect 7573 12189 7607 12223
rect 8125 12189 8159 12223
rect 8217 12189 8251 12223
rect 8677 12189 8711 12223
rect 10333 12189 10367 12223
rect 10426 12189 10460 12223
rect 10839 12189 10873 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 11345 12199 11379 12233
rect 11529 12189 11563 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12081 12189 12115 12223
rect 12173 12189 12207 12223
rect 13921 12189 13955 12223
rect 2145 12121 2179 12155
rect 2237 12121 2271 12155
rect 4245 12121 4279 12155
rect 4445 12121 4479 12155
rect 4997 12121 5031 12155
rect 5917 12121 5951 12155
rect 7849 12121 7883 12155
rect 8401 12121 8435 12155
rect 9597 12121 9631 12155
rect 10609 12121 10643 12155
rect 10701 12121 10735 12155
rect 11161 12121 11195 12155
rect 13277 12121 13311 12155
rect 13461 12121 13495 12155
rect 13829 12121 13863 12155
rect 2697 12053 2731 12087
rect 4077 12053 4111 12087
rect 4629 12053 4663 12087
rect 4797 12053 4831 12087
rect 5641 12053 5675 12087
rect 5825 12053 5859 12087
rect 6009 12053 6043 12087
rect 6653 12053 6687 12087
rect 7941 12053 7975 12087
rect 8585 12053 8619 12087
rect 10057 12053 10091 12087
rect 4537 11849 4571 11883
rect 4705 11849 4739 11883
rect 4997 11849 5031 11883
rect 5165 11849 5199 11883
rect 5625 11849 5659 11883
rect 13461 11849 13495 11883
rect 4905 11781 4939 11815
rect 5365 11781 5399 11815
rect 5825 11781 5859 11815
rect 10793 11781 10827 11815
rect 13553 11781 13587 11815
rect 3985 11713 4019 11747
rect 8585 11713 8619 11747
rect 10701 11713 10735 11747
rect 11069 11713 11103 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 11621 11713 11655 11747
rect 11897 11713 11931 11747
rect 12265 11713 12299 11747
rect 12449 11713 12483 11747
rect 12541 11713 12575 11747
rect 12817 11713 12851 11747
rect 3801 11645 3835 11679
rect 11713 11645 11747 11679
rect 12633 11645 12667 11679
rect 13185 11645 13219 11679
rect 5457 11577 5491 11611
rect 11897 11577 11931 11611
rect 13001 11577 13035 11611
rect 13277 11577 13311 11611
rect 4169 11509 4203 11543
rect 4721 11509 4755 11543
rect 5181 11509 5215 11543
rect 5641 11509 5675 11543
rect 8769 11509 8803 11543
rect 13093 11509 13127 11543
rect 3801 11305 3835 11339
rect 8309 11305 8343 11339
rect 8769 11305 8803 11339
rect 9413 11305 9447 11339
rect 1961 11237 1995 11271
rect 2329 11237 2363 11271
rect 7481 11237 7515 11271
rect 7757 11237 7791 11271
rect 9045 11237 9079 11271
rect 1777 11169 1811 11203
rect 2513 11169 2547 11203
rect 4445 11169 4479 11203
rect 6285 11169 6319 11203
rect 7849 11169 7883 11203
rect 8677 11169 8711 11203
rect 2605 11101 2639 11135
rect 2697 11101 2731 11135
rect 2789 11101 2823 11135
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 4537 11101 4571 11135
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5273 11101 5307 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6193 11101 6227 11135
rect 6561 11101 6595 11135
rect 6653 11101 6687 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 7941 11101 7975 11135
rect 8217 11101 8251 11135
rect 8493 11101 8527 11135
rect 9229 11101 9263 11135
rect 9689 11101 9723 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 10057 11101 10091 11135
rect 2237 11033 2271 11067
rect 8769 11033 8803 11067
rect 10793 11033 10827 11067
rect 4169 10965 4203 10999
rect 4629 10965 4663 10999
rect 5457 10965 5491 10999
rect 8125 10965 8159 10999
rect 12265 10965 12299 10999
rect 2145 10761 2179 10795
rect 2605 10761 2639 10795
rect 2697 10761 2731 10795
rect 3985 10761 4019 10795
rect 5273 10761 5307 10795
rect 6469 10761 6503 10795
rect 9045 10761 9079 10795
rect 9597 10761 9631 10795
rect 10425 10761 10459 10795
rect 11177 10761 11211 10795
rect 11345 10761 11379 10795
rect 13921 10761 13955 10795
rect 5089 10693 5123 10727
rect 5365 10693 5399 10727
rect 9413 10693 9447 10727
rect 10977 10693 11011 10727
rect 12808 10693 12842 10727
rect 2329 10625 2363 10659
rect 2789 10625 2823 10659
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 3893 10625 3927 10659
rect 4169 10625 4203 10659
rect 5457 10625 5491 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 8677 10625 8711 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 9781 10625 9815 10659
rect 10241 10625 10275 10659
rect 10333 10625 10367 10659
rect 10609 10625 10643 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 2421 10557 2455 10591
rect 4261 10557 4295 10591
rect 8769 10557 8803 10591
rect 9965 10557 9999 10591
rect 11529 10557 11563 10591
rect 12541 10557 12575 10591
rect 5641 10489 5675 10523
rect 11805 10489 11839 10523
rect 8861 10421 8895 10455
rect 9965 10421 9999 10455
rect 10609 10421 10643 10455
rect 11161 10421 11195 10455
rect 4445 10217 4479 10251
rect 6837 10217 6871 10251
rect 7573 10217 7607 10251
rect 10885 10217 10919 10251
rect 13737 10217 13771 10251
rect 2789 10149 2823 10183
rect 7757 10149 7791 10183
rect 4629 10081 4663 10115
rect 6745 10081 6779 10115
rect 6929 10081 6963 10115
rect 7481 10081 7515 10115
rect 1409 10013 1443 10047
rect 4077 10013 4111 10047
rect 4537 10013 4571 10047
rect 7205 10013 7239 10047
rect 7297 10013 7331 10047
rect 7573 10013 7607 10047
rect 8217 10013 8251 10047
rect 10885 10013 10919 10047
rect 11161 10013 11195 10047
rect 12173 10013 12207 10047
rect 12357 10013 12391 10047
rect 1676 9945 1710 9979
rect 4169 9945 4203 9979
rect 6377 9945 6411 9979
rect 8309 9945 8343 9979
rect 12817 9945 12851 9979
rect 13185 9945 13219 9979
rect 13369 9945 13403 9979
rect 13553 9945 13587 9979
rect 3801 9877 3835 9911
rect 4261 9877 4295 9911
rect 6469 9877 6503 9911
rect 7113 9877 7147 9911
rect 11069 9877 11103 9911
rect 12265 9877 12299 9911
rect 1777 9673 1811 9707
rect 4997 9673 5031 9707
rect 7389 9673 7423 9707
rect 11805 9673 11839 9707
rect 4905 9605 4939 9639
rect 5365 9605 5399 9639
rect 6929 9605 6963 9639
rect 10425 9605 10459 9639
rect 1961 9537 1995 9571
rect 3157 9537 3191 9571
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 5762 9537 5796 9571
rect 6101 9537 6135 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 7849 9537 7883 9571
rect 8769 9537 8803 9571
rect 9321 9537 9355 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11529 9537 11563 9571
rect 12081 9537 12115 9571
rect 12265 9537 12299 9571
rect 12357 9537 12391 9571
rect 12449 9537 12483 9571
rect 12817 9537 12851 9571
rect 13073 9537 13107 9571
rect 3249 9469 3283 9503
rect 3341 9469 3375 9503
rect 3433 9469 3467 9503
rect 4629 9469 4663 9503
rect 5114 9469 5148 9503
rect 9045 9469 9079 9503
rect 11805 9469 11839 9503
rect 4261 9401 4295 9435
rect 4353 9401 4387 9435
rect 5273 9401 5307 9435
rect 5963 9401 5997 9435
rect 12725 9401 12759 9435
rect 2973 9333 3007 9367
rect 5825 9333 5859 9367
rect 6469 9333 6503 9367
rect 6653 9333 6687 9367
rect 8309 9333 8343 9367
rect 8953 9333 8987 9367
rect 11621 9333 11655 9367
rect 14197 9333 14231 9367
rect 6101 9129 6135 9163
rect 2421 9061 2455 9095
rect 8769 9061 8803 9095
rect 11253 9061 11287 9095
rect 11529 9061 11563 9095
rect 12357 9061 12391 9095
rect 2881 8993 2915 9027
rect 3249 8993 3283 9027
rect 3893 8993 3927 9027
rect 6469 8993 6503 9027
rect 9321 8993 9355 9027
rect 9413 8993 9447 9027
rect 9873 8993 9907 9027
rect 2789 8925 2823 8959
rect 3157 8925 3191 8959
rect 4169 8925 4203 8959
rect 4537 8925 4571 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 7021 8925 7055 8959
rect 7297 8925 7331 8959
rect 7481 8925 7515 8959
rect 8125 8925 8159 8959
rect 8217 8925 8251 8959
rect 8585 8925 8619 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 9597 8925 9631 8959
rect 11345 8925 11379 8959
rect 12357 8925 12391 8959
rect 12817 8925 12851 8959
rect 13093 8925 13127 8959
rect 2053 8857 2087 8891
rect 2605 8857 2639 8891
rect 5733 8857 5767 8891
rect 5917 8857 5951 8891
rect 8401 8857 8435 8891
rect 8493 8857 8527 8891
rect 9781 8857 9815 8891
rect 10118 8857 10152 8891
rect 2513 8789 2547 8823
rect 3065 8789 3099 8823
rect 6837 8789 6871 8823
rect 7205 8789 7239 8823
rect 10057 8585 10091 8619
rect 12173 8585 12207 8619
rect 2513 8449 2547 8483
rect 5733 8449 5767 8483
rect 5825 8449 5859 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 12725 8449 12759 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 7849 8381 7883 8415
rect 2329 8245 2363 8279
rect 5457 8245 5491 8279
rect 5825 8245 5859 8279
rect 6561 8245 6595 8279
rect 9689 8245 9723 8279
rect 4169 8041 4203 8075
rect 4629 8041 4663 8075
rect 6653 8041 6687 8075
rect 7297 8041 7331 8075
rect 8677 8041 8711 8075
rect 9321 8041 9355 8075
rect 10333 8041 10367 8075
rect 8953 7973 8987 8007
rect 11069 7973 11103 8007
rect 2053 7905 2087 7939
rect 5340 7905 5374 7939
rect 6837 7905 6871 7939
rect 7389 7905 7423 7939
rect 3801 7837 3835 7871
rect 3893 7837 3927 7871
rect 4261 7837 4295 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6193 7837 6227 7871
rect 6377 7837 6411 7871
rect 6469 7837 6503 7871
rect 6561 7837 6595 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 8401 7837 8435 7871
rect 9413 7837 9447 7871
rect 10241 7837 10275 7871
rect 10333 7837 10367 7871
rect 10609 7837 10643 7871
rect 11161 7837 11195 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 2320 7769 2354 7803
rect 5457 7769 5491 7803
rect 6837 7769 6871 7803
rect 8677 7769 8711 7803
rect 9873 7769 9907 7803
rect 3433 7701 3467 7735
rect 3985 7701 4019 7735
rect 4261 7701 4295 7735
rect 5181 7701 5215 7735
rect 5549 7701 5583 7735
rect 7021 7701 7055 7735
rect 7665 7701 7699 7735
rect 8493 7701 8527 7735
rect 10517 7701 10551 7735
rect 3623 7497 3657 7531
rect 5365 7497 5399 7531
rect 3709 7429 3743 7463
rect 6101 7429 6135 7463
rect 7481 7429 7515 7463
rect 11529 7429 11563 7463
rect 3525 7361 3559 7395
rect 3801 7351 3835 7385
rect 5273 7361 5307 7395
rect 5457 7361 5491 7395
rect 8309 7361 8343 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 9137 7361 9171 7395
rect 9597 7361 9631 7395
rect 9689 7361 9723 7395
rect 10609 7361 10643 7395
rect 7849 7293 7883 7327
rect 8401 7293 8435 7327
rect 9873 7293 9907 7327
rect 8769 7225 8803 7259
rect 5825 7157 5859 7191
rect 7941 7157 7975 7191
rect 9781 7157 9815 7191
rect 10425 7157 10459 7191
rect 12817 7157 12851 7191
rect 5181 6953 5215 6987
rect 7297 6953 7331 6987
rect 10149 6953 10183 6987
rect 7665 6885 7699 6919
rect 10241 6885 10275 6919
rect 3801 6817 3835 6851
rect 5621 6817 5655 6851
rect 9597 6817 9631 6851
rect 9781 6817 9815 6851
rect 10057 6817 10091 6851
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 6173 6749 6207 6783
rect 7665 6749 7699 6783
rect 7941 6749 7975 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 9459 6749 9493 6783
rect 10609 6749 10643 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 4068 6681 4102 6715
rect 5549 6681 5583 6715
rect 9229 6681 9263 6715
rect 11774 6681 11808 6715
rect 5365 6613 5399 6647
rect 8953 6613 8987 6647
rect 11253 6613 11287 6647
rect 12909 6613 12943 6647
rect 8493 6409 8527 6443
rect 11062 6409 11096 6443
rect 2228 6341 2262 6375
rect 8033 6341 8067 6375
rect 8677 6341 8711 6375
rect 3617 6273 3651 6307
rect 4905 6273 4939 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 5825 6273 5859 6307
rect 7849 6273 7883 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8769 6273 8803 6307
rect 9781 6273 9815 6307
rect 9959 6273 9993 6307
rect 10045 6283 10079 6317
rect 10241 6273 10275 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11713 6283 11747 6317
rect 11897 6273 11931 6307
rect 12265 6273 12299 6307
rect 13665 6273 13699 6307
rect 13921 6273 13955 6307
rect 1961 6205 1995 6239
rect 3801 6205 3835 6239
rect 5181 6205 5215 6239
rect 5365 6205 5399 6239
rect 10333 6205 10367 6239
rect 10425 6205 10459 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 12449 6205 12483 6239
rect 9781 6137 9815 6171
rect 3341 6069 3375 6103
rect 3433 6069 3467 6103
rect 6009 6069 6043 6103
rect 7665 6069 7699 6103
rect 10793 6069 10827 6103
rect 12541 6069 12575 6103
rect 2421 5865 2455 5899
rect 3801 5865 3835 5899
rect 4997 5865 5031 5899
rect 8217 5865 8251 5899
rect 8677 5865 8711 5899
rect 9321 5865 9355 5899
rect 11621 5865 11655 5899
rect 12357 5865 12391 5899
rect 11713 5797 11747 5831
rect 12173 5797 12207 5831
rect 9413 5729 9447 5763
rect 10149 5729 10183 5763
rect 11805 5729 11839 5763
rect 2605 5661 2639 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 4353 5661 4387 5695
rect 4445 5661 4479 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 6837 5661 6871 5695
rect 7205 5661 7239 5695
rect 7665 5661 7699 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 9321 5661 9355 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 11253 5661 11287 5695
rect 11437 5661 11471 5695
rect 11529 5661 11563 5695
rect 12541 5661 12575 5695
rect 12808 5661 12842 5695
rect 4169 5593 4203 5627
rect 4629 5593 4663 5627
rect 6929 5593 6963 5627
rect 7849 5593 7883 5627
rect 9873 5593 9907 5627
rect 10333 5593 10367 5627
rect 11897 5593 11931 5627
rect 5549 5525 5583 5559
rect 9689 5525 9723 5559
rect 11345 5525 11379 5559
rect 13921 5525 13955 5559
rect 3801 5321 3835 5355
rect 4813 5321 4847 5355
rect 9045 5321 9079 5355
rect 13645 5321 13679 5355
rect 3525 5253 3559 5287
rect 3249 5185 3283 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 5937 5185 5971 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 7665 5185 7699 5219
rect 8953 5185 8987 5219
rect 9137 5185 9171 5219
rect 10701 5185 10735 5219
rect 10885 5185 10919 5219
rect 11897 5185 11931 5219
rect 12173 5185 12207 5219
rect 12909 5185 12943 5219
rect 13185 5185 13219 5219
rect 13553 5185 13587 5219
rect 13829 5185 13863 5219
rect 4261 5117 4295 5151
rect 6193 5117 6227 5151
rect 7941 5117 7975 5151
rect 12725 5117 12759 5151
rect 6469 5049 6503 5083
rect 3893 4981 3927 5015
rect 7849 4981 7883 5015
rect 8217 4981 8251 5015
rect 10701 4981 10735 5015
rect 11989 4981 12023 5015
rect 12449 4981 12483 5015
rect 14013 4981 14047 5015
rect 11805 4777 11839 4811
rect 12265 4777 12299 4811
rect 9137 4709 9171 4743
rect 1593 4573 1627 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 6469 4573 6503 4607
rect 6745 4573 6779 4607
rect 6837 4573 6871 4607
rect 9229 4573 9263 4607
rect 10425 4573 10459 4607
rect 12541 4573 12575 4607
rect 1860 4505 1894 4539
rect 4169 4505 4203 4539
rect 6653 4505 6687 4539
rect 8953 4505 8987 4539
rect 10670 4505 10704 4539
rect 12081 4505 12115 4539
rect 12297 4505 12331 4539
rect 12808 4505 12842 4539
rect 2973 4437 3007 4471
rect 3801 4437 3835 4471
rect 7021 4437 7055 4471
rect 9229 4437 9263 4471
rect 12449 4437 12483 4471
rect 13921 4437 13955 4471
rect 2053 4233 2087 4267
rect 5457 4233 5491 4267
rect 8309 4233 8343 4267
rect 8953 4233 8987 4267
rect 12817 4233 12851 4267
rect 13645 4233 13679 4267
rect 4445 4165 4479 4199
rect 5089 4165 5123 4199
rect 5181 4165 5215 4199
rect 6745 4165 6779 4199
rect 8401 4165 8435 4199
rect 9873 4165 9907 4199
rect 2237 4097 2271 4131
rect 3433 4097 3467 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 4629 4097 4663 4131
rect 4905 4097 4939 4131
rect 5273 4097 5307 4131
rect 5733 4097 5767 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 8125 4097 8159 4131
rect 9045 4097 9079 4131
rect 9321 4097 9355 4131
rect 9597 4097 9631 4131
rect 9778 4119 9812 4153
rect 10057 4097 10091 4131
rect 10793 4097 10827 4131
rect 12633 4097 12667 4131
rect 13553 4097 13587 4131
rect 3617 4029 3651 4063
rect 5917 4029 5951 4063
rect 7021 4029 7055 4063
rect 8033 4029 8067 4063
rect 9413 4029 9447 4063
rect 10517 4029 10551 4063
rect 10977 4029 11011 4063
rect 9505 3961 9539 3995
rect 3249 3893 3283 3927
rect 4813 3893 4847 3927
rect 5549 3893 5583 3927
rect 6377 3893 6411 3927
rect 7389 3893 7423 3927
rect 7941 3893 7975 3927
rect 9137 3893 9171 3927
rect 10241 3893 10275 3927
rect 10609 3893 10643 3927
rect 9781 3689 9815 3723
rect 5549 3553 5583 3587
rect 2881 3485 2915 3519
rect 4629 3485 4663 3519
rect 4813 3485 4847 3519
rect 5733 3485 5767 3519
rect 6009 3485 6043 3519
rect 7665 3485 7699 3519
rect 9505 3485 9539 3519
rect 9597 3485 9631 3519
rect 6276 3417 6310 3451
rect 9781 3417 9815 3451
rect 2697 3349 2731 3383
rect 4445 3349 4479 3383
rect 5917 3349 5951 3383
rect 7389 3349 7423 3383
rect 7481 3349 7515 3383
rect 4537 3145 4571 3179
rect 6009 3145 6043 3179
rect 6377 3145 6411 3179
rect 9137 3145 9171 3179
rect 10425 3145 10459 3179
rect 14013 3145 14047 3179
rect 8002 3077 8036 3111
rect 3157 3009 3191 3043
rect 3424 3009 3458 3043
rect 4629 3009 4663 3043
rect 4896 3009 4930 3043
rect 6561 3009 6595 3043
rect 7757 3009 7791 3043
rect 10701 3009 10735 3043
rect 12633 3009 12667 3043
rect 12900 3009 12934 3043
rect 10885 2805 10919 2839
rect 3801 2601 3835 2635
rect 4997 2601 5031 2635
rect 8585 2601 8619 2635
rect 10609 2601 10643 2635
rect 13461 2601 13495 2635
rect 3617 2533 3651 2567
rect 2237 2465 2271 2499
rect 7205 2465 7239 2499
rect 1593 2397 1627 2431
rect 2145 2397 2179 2431
rect 2504 2397 2538 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 6193 2397 6227 2431
rect 6929 2397 6963 2431
rect 7472 2397 7506 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 10885 2397 10919 2431
rect 11345 2397 11379 2431
rect 12633 2397 12667 2431
rect 13645 2397 13679 2431
rect 13921 2397 13955 2431
rect 9474 2329 9508 2363
rect 1409 2261 1443 2295
rect 1961 2261 1995 2295
rect 4077 2261 4111 2295
rect 4721 2261 4755 2295
rect 6009 2261 6043 2295
rect 7113 2261 7147 2295
rect 8953 2261 8987 2295
rect 10701 2261 10735 2295
rect 11161 2261 11195 2295
rect 12449 2261 12483 2295
rect 13737 2261 13771 2295
<< metal1 >>
rect 1104 15258 14536 15280
rect 1104 15206 4918 15258
rect 4970 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 5238 15258
rect 5290 15206 10918 15258
rect 10970 15206 10982 15258
rect 11034 15206 11046 15258
rect 11098 15206 11110 15258
rect 11162 15206 11174 15258
rect 11226 15206 11238 15258
rect 11290 15206 14536 15258
rect 1104 15184 14536 15206
rect 658 15104 664 15156
rect 716 15144 722 15156
rect 1397 15147 1455 15153
rect 1397 15144 1409 15147
rect 716 15116 1409 15144
rect 716 15104 722 15116
rect 1397 15113 1409 15116
rect 1443 15113 1455 15147
rect 1397 15107 1455 15113
rect 1854 15104 1860 15156
rect 1912 15104 1918 15156
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2924 15116 2973 15144
rect 2924 15104 2930 15116
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 4028 15116 4077 15144
rect 4028 15104 4034 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 5169 15147 5227 15153
rect 5169 15113 5181 15147
rect 5215 15144 5227 15147
rect 5350 15144 5356 15156
rect 5215 15116 5356 15144
rect 5215 15113 5227 15116
rect 5169 15107 5227 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 6236 15116 6377 15144
rect 6236 15104 6242 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 7374 15104 7380 15156
rect 7432 15104 7438 15156
rect 8478 15104 8484 15156
rect 8536 15104 8542 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 9548 15116 9597 15144
rect 9548 15104 9554 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 11698 15104 11704 15156
rect 11756 15104 11762 15156
rect 12802 15104 12808 15156
rect 12860 15104 12866 15156
rect 3602 15076 3608 15088
rect 2056 15048 3608 15076
rect 1578 14968 1584 15020
rect 1636 14968 1642 15020
rect 2056 15017 2084 15048
rect 3602 15036 3608 15048
rect 3660 15036 3666 15088
rect 4706 15036 4712 15088
rect 4764 15076 4770 15088
rect 4764 15048 7604 15076
rect 4764 15036 4770 15048
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 3418 15008 3424 15020
rect 3191 14980 3424 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 4246 14968 4252 15020
rect 4304 14968 4310 15020
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 7576 15017 7604 15048
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 4396 14980 5365 15008
rect 4396 14968 4402 14980
rect 5353 14977 5365 14980
rect 5399 14977 5411 15011
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5353 14971 5411 14977
rect 5460 14980 6561 15008
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 5460 14940 5488 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 14977 7619 15011
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 7561 14971 7619 14977
rect 7668 14980 8677 15008
rect 3292 14912 5488 14940
rect 3292 14900 3298 14912
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 7668 14940 7696 14980
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 6696 14912 7696 14940
rect 6696 14900 6702 14912
rect 7834 14900 7840 14952
rect 7892 14940 7898 14952
rect 9784 14940 9812 14971
rect 7892 14912 9812 14940
rect 10336 14940 10364 14971
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 11716 15008 11744 15104
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11716 14980 11805 15008
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 12820 15008 12848 15104
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 12820 14980 12909 15008
rect 11793 14971 11851 14977
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 13906 14968 13912 15020
rect 13964 14968 13970 15020
rect 10336 14912 12940 14940
rect 7892 14900 7898 14912
rect 5442 14832 5448 14884
rect 5500 14872 5506 14884
rect 10336 14872 10364 14912
rect 5500 14844 10364 14872
rect 5500 14832 5506 14844
rect 12912 14816 12940 14912
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 10686 14804 10692 14816
rect 10551 14776 10692 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11974 14764 11980 14816
rect 12032 14764 12038 14816
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13078 14764 13084 14816
rect 13136 14764 13142 14816
rect 13722 14764 13728 14816
rect 13780 14764 13786 14816
rect 1104 14714 14536 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13918 14714
rect 13970 14662 13982 14714
rect 14034 14662 14046 14714
rect 14098 14662 14110 14714
rect 14162 14662 14174 14714
rect 14226 14662 14238 14714
rect 14290 14662 14536 14714
rect 1104 14640 14536 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 1636 14572 7389 14600
rect 1636 14560 1642 14572
rect 7377 14569 7389 14572
rect 7423 14600 7435 14603
rect 8938 14600 8944 14612
rect 7423 14572 8944 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 13722 14600 13728 14612
rect 9272 14572 13728 14600
rect 9272 14560 9278 14572
rect 3234 14492 3240 14544
rect 3292 14492 3298 14544
rect 12176 14436 12388 14464
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1544 14368 1869 14396
rect 1544 14356 1550 14368
rect 1857 14365 1869 14368
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 3510 14356 3516 14408
rect 3568 14396 3574 14408
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 3568 14368 5181 14396
rect 3568 14356 3574 14368
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9033 14399 9091 14405
rect 9033 14396 9045 14399
rect 8812 14368 9045 14396
rect 8812 14356 8818 14368
rect 9033 14365 9045 14368
rect 9079 14365 9091 14399
rect 9033 14359 9091 14365
rect 9300 14399 9358 14405
rect 9300 14365 9312 14399
rect 9346 14396 9358 14399
rect 10597 14399 10655 14405
rect 9346 14368 9536 14396
rect 9346 14365 9358 14368
rect 9300 14359 9358 14365
rect 2124 14331 2182 14337
rect 2124 14297 2136 14331
rect 2170 14328 2182 14331
rect 2222 14328 2228 14340
rect 2170 14300 2228 14328
rect 2170 14297 2182 14300
rect 2124 14291 2182 14297
rect 2222 14288 2228 14300
rect 2280 14288 2286 14340
rect 5436 14331 5494 14337
rect 5436 14297 5448 14331
rect 5482 14328 5494 14331
rect 5626 14328 5632 14340
rect 5482 14300 5632 14328
rect 5482 14297 5494 14300
rect 5436 14291 5494 14297
rect 5626 14288 5632 14300
rect 5684 14288 5690 14340
rect 8478 14288 8484 14340
rect 8536 14337 8542 14340
rect 8536 14291 8548 14337
rect 8536 14288 8542 14291
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 4856 14232 6561 14260
rect 4856 14220 4862 14232
rect 6549 14229 6561 14232
rect 6595 14260 6607 14263
rect 6638 14260 6644 14272
rect 6595 14232 6644 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 9048 14260 9076 14359
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9508 14328 9536 14368
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10643 14368 11008 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10612 14328 10640 14359
rect 9456 14300 9536 14328
rect 9600 14300 10640 14328
rect 9456 14288 9462 14300
rect 9600 14260 9628 14300
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 10842 14331 10900 14337
rect 10842 14328 10854 14331
rect 10744 14300 10854 14328
rect 10744 14288 10750 14300
rect 10842 14297 10854 14300
rect 10888 14297 10900 14331
rect 10980 14328 11008 14368
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 12176 14396 12204 14436
rect 11480 14368 12204 14396
rect 11480 14356 11486 14368
rect 12250 14356 12256 14408
rect 12308 14356 12314 14408
rect 12360 14396 12388 14436
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 12360 14368 12541 14396
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12710 14356 12716 14408
rect 12768 14356 12774 14408
rect 12912 14405 12940 14572
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 12728 14328 12756 14356
rect 10980 14300 12756 14328
rect 10842 14291 10900 14297
rect 9048 14232 9628 14260
rect 10410 14220 10416 14272
rect 10468 14220 10474 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11848 14232 11989 14260
rect 11848 14220 11854 14232
rect 11977 14229 11989 14232
rect 12023 14260 12035 14263
rect 12066 14260 12072 14272
rect 12023 14232 12072 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12158 14220 12164 14272
rect 12216 14260 12222 14272
rect 12342 14260 12348 14272
rect 12216 14232 12348 14260
rect 12216 14220 12222 14232
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 12676 14232 12725 14260
rect 12676 14220 12682 14232
rect 12713 14229 12725 14232
rect 12759 14229 12771 14263
rect 12713 14223 12771 14229
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12952 14232 13001 14260
rect 12952 14220 12958 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 12989 14223 13047 14229
rect 1104 14170 14536 14192
rect 1104 14118 4918 14170
rect 4970 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 5238 14170
rect 5290 14118 10918 14170
rect 10970 14118 10982 14170
rect 11034 14118 11046 14170
rect 11098 14118 11110 14170
rect 11162 14118 11174 14170
rect 11226 14118 11238 14170
rect 11290 14118 14536 14170
rect 1104 14096 14536 14118
rect 2222 14016 2228 14068
rect 2280 14016 2286 14068
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 2547 14028 3157 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 3145 14025 3157 14028
rect 3191 14025 3203 14059
rect 3145 14019 3203 14025
rect 3421 14059 3479 14065
rect 3421 14025 3433 14059
rect 3467 14056 3479 14059
rect 3467 14028 3832 14056
rect 3467 14025 3479 14028
rect 3421 14019 3479 14025
rect 2516 13932 2544 14019
rect 2593 13991 2651 13997
rect 2593 13957 2605 13991
rect 2639 13988 2651 13991
rect 3694 13988 3700 14000
rect 2639 13960 3096 13988
rect 2639 13957 2651 13960
rect 2593 13951 2651 13957
rect 3068 13932 3096 13960
rect 3436 13960 3700 13988
rect 2222 13880 2228 13932
rect 2280 13880 2286 13932
rect 2498 13880 2504 13932
rect 2556 13880 2562 13932
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2866 13920 2872 13932
rect 2731 13892 2872 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 2958 13880 2964 13932
rect 3016 13880 3022 13932
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 3436 13929 3464 13960
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 3804 13988 3832 14028
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4764 14028 4997 14056
rect 4764 14016 4770 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 6089 14059 6147 14065
rect 6089 14056 6101 14059
rect 5316 14028 6101 14056
rect 5316 14016 5322 14028
rect 6089 14025 6101 14028
rect 6135 14025 6147 14059
rect 6089 14019 6147 14025
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7892 14028 8033 14056
rect 7892 14016 7898 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8536 14028 8585 14056
rect 8536 14016 8542 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 8573 14019 8631 14025
rect 10502 14016 10508 14068
rect 10560 14016 10566 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 12158 14016 12164 14068
rect 12216 14016 12222 14068
rect 12443 14059 12501 14065
rect 12443 14025 12455 14059
rect 12489 14025 12501 14059
rect 12443 14019 12501 14025
rect 12529 14059 12587 14065
rect 12529 14025 12541 14059
rect 12575 14056 12587 14059
rect 12618 14056 12624 14068
rect 12575 14028 12624 14056
rect 12575 14025 12587 14028
rect 12529 14019 12587 14025
rect 3861 13991 3919 13997
rect 3861 13988 3873 13991
rect 3804 13960 3873 13988
rect 3861 13957 3873 13960
rect 3907 13957 3919 13991
rect 9858 13988 9864 14000
rect 3861 13951 3919 13957
rect 4080 13960 6684 13988
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 4080 13920 4108 13960
rect 3421 13883 3479 13889
rect 3620 13892 4108 13920
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 3510 13852 3516 13864
rect 1544 13824 3516 13852
rect 1544 13812 1550 13824
rect 3510 13812 3516 13824
rect 3568 13852 3574 13864
rect 3620 13861 3648 13892
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4798 13920 4804 13932
rect 4212 13892 4804 13920
rect 4212 13880 4218 13892
rect 4798 13880 4804 13892
rect 4856 13920 4862 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4856 13892 5089 13920
rect 4856 13880 4862 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5258 13880 5264 13932
rect 5316 13880 5322 13932
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5721 13928 5779 13929
rect 5644 13923 5779 13928
rect 5644 13920 5733 13923
rect 5500 13900 5733 13920
rect 5500 13892 5672 13900
rect 5500 13880 5506 13892
rect 3605 13855 3663 13861
rect 3605 13852 3617 13855
rect 3568 13824 3617 13852
rect 3568 13812 3574 13824
rect 3605 13821 3617 13824
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 3016 13756 3464 13784
rect 3016 13744 3022 13756
rect 2317 13719 2375 13725
rect 2317 13685 2329 13719
rect 2363 13716 2375 13719
rect 3142 13716 3148 13728
rect 2363 13688 3148 13716
rect 2363 13685 2375 13688
rect 2317 13679 2375 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3326 13676 3332 13728
rect 3384 13676 3390 13728
rect 3436 13716 3464 13756
rect 4982 13744 4988 13796
rect 5040 13784 5046 13796
rect 5552 13784 5580 13892
rect 5721 13889 5733 13900
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 5810 13880 5816 13932
rect 5868 13920 5874 13932
rect 5951 13923 6009 13929
rect 5951 13920 5963 13923
rect 5868 13892 5963 13920
rect 5868 13880 5874 13892
rect 5951 13889 5963 13892
rect 5997 13889 6009 13923
rect 5951 13883 6009 13889
rect 6178 13880 6184 13932
rect 6236 13880 6242 13932
rect 6656 13929 6684 13960
rect 8864 13960 9864 13988
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6897 13923 6955 13929
rect 6897 13920 6909 13923
rect 6641 13883 6699 13889
rect 6748 13892 6909 13920
rect 6748 13852 6776 13892
rect 6897 13889 6909 13892
rect 6943 13889 6955 13923
rect 6897 13883 6955 13889
rect 8864 13861 8892 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 11808 13988 11836 14016
rect 12176 13988 12204 14016
rect 11716 13960 11836 13988
rect 11992 13960 12204 13988
rect 12452 13988 12480 14019
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12958 13991 13016 13997
rect 12958 13988 12970 13991
rect 12452 13960 12970 13988
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9309 13923 9367 13929
rect 9309 13920 9321 13923
rect 9272 13892 9321 13920
rect 9272 13880 9278 13892
rect 9309 13889 9321 13892
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9950 13920 9956 13932
rect 9539 13892 9956 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10686 13923 10744 13929
rect 10686 13889 10698 13923
rect 10732 13920 10744 13923
rect 11330 13920 11336 13932
rect 10732 13892 11336 13920
rect 10732 13889 10744 13892
rect 10686 13883 10744 13889
rect 11330 13880 11336 13892
rect 11388 13920 11394 13932
rect 11716 13929 11744 13960
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11388 13892 11713 13920
rect 11388 13880 11394 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 11992 13929 12020 13960
rect 12958 13957 12970 13960
rect 13004 13957 13016 13991
rect 12958 13951 13016 13957
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 11848 13892 11897 13920
rect 11848 13880 11854 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12335 13923 12393 13929
rect 12335 13920 12347 13923
rect 12268 13892 12347 13920
rect 5828 13824 6776 13852
rect 8757 13855 8815 13861
rect 5040 13756 5580 13784
rect 5721 13787 5779 13793
rect 5040 13744 5046 13756
rect 5721 13753 5733 13787
rect 5767 13784 5779 13787
rect 5828 13784 5856 13824
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9398 13852 9404 13864
rect 9079 13824 9404 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 5767 13756 5856 13784
rect 8772 13784 8800 13815
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 10134 13812 10140 13864
rect 10192 13852 10198 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 10192 13824 11161 13852
rect 10192 13812 10198 13824
rect 11149 13821 11161 13824
rect 11195 13852 11207 13855
rect 11422 13852 11428 13864
rect 11195 13824 11428 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 11698 13784 11704 13796
rect 8772 13756 11704 13784
rect 5767 13753 5779 13756
rect 5721 13747 5779 13753
rect 11698 13744 11704 13756
rect 11756 13784 11762 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11756 13756 11805 13784
rect 11756 13744 11762 13756
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 3878 13716 3884 13728
rect 3436 13688 3884 13716
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 5000 13716 5028 13744
rect 4028 13688 5028 13716
rect 4028 13676 4034 13688
rect 5074 13676 5080 13728
rect 5132 13676 5138 13728
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5626 13716 5632 13728
rect 5224 13688 5632 13716
rect 5224 13676 5230 13688
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 5813 13719 5871 13725
rect 5813 13685 5825 13719
rect 5859 13716 5871 13719
rect 6546 13716 6552 13728
rect 5859 13688 6552 13716
rect 5859 13685 5871 13688
rect 5813 13679 5871 13685
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13716 11115 13719
rect 11517 13719 11575 13725
rect 11517 13716 11529 13719
rect 11103 13688 11529 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 11517 13685 11529 13688
rect 11563 13685 11575 13719
rect 12268 13716 12296 13892
rect 12335 13889 12347 13892
rect 12381 13889 12393 13923
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12335 13883 12393 13889
rect 12544 13892 12633 13920
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12544 13852 12572 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 12492 13824 12572 13852
rect 12492 13812 12498 13824
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 12894 13716 12900 13728
rect 12268 13688 12900 13716
rect 11517 13679 11575 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14093 13719 14151 13725
rect 14093 13716 14105 13719
rect 13872 13688 14105 13716
rect 13872 13676 13878 13688
rect 14093 13685 14105 13688
rect 14139 13685 14151 13719
rect 14093 13679 14151 13685
rect 1104 13626 14536 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13918 13626
rect 13970 13574 13982 13626
rect 14034 13574 14046 13626
rect 14098 13574 14110 13626
rect 14162 13574 14174 13626
rect 14226 13574 14238 13626
rect 14290 13574 14536 13626
rect 1104 13552 14536 13574
rect 3142 13472 3148 13524
rect 3200 13472 3206 13524
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3384 13484 4077 13512
rect 3384 13472 3390 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4985 13515 5043 13521
rect 4985 13481 4997 13515
rect 5031 13512 5043 13515
rect 5074 13512 5080 13524
rect 5031 13484 5080 13512
rect 5031 13481 5043 13484
rect 4985 13475 5043 13481
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 6546 13472 6552 13524
rect 6604 13472 6610 13524
rect 7834 13472 7840 13524
rect 7892 13472 7898 13524
rect 9585 13515 9643 13521
rect 9585 13481 9597 13515
rect 9631 13512 9643 13515
rect 9674 13512 9680 13524
rect 9631 13484 9680 13512
rect 9631 13481 9643 13484
rect 9585 13475 9643 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 11698 13512 11704 13524
rect 11480 13484 11704 13512
rect 11480 13472 11486 13484
rect 11698 13472 11704 13484
rect 11756 13512 11762 13524
rect 11793 13515 11851 13521
rect 11793 13512 11805 13515
rect 11756 13484 11805 13512
rect 11756 13472 11762 13484
rect 11793 13481 11805 13484
rect 11839 13481 11851 13515
rect 11793 13475 11851 13481
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 2498 13404 2504 13456
rect 2556 13444 2562 13456
rect 4893 13447 4951 13453
rect 2556 13416 4660 13444
rect 2556 13404 2562 13416
rect 4338 13376 4344 13388
rect 2792 13348 4344 13376
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1486 13308 1492 13320
rect 1443 13280 1492 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 1670 13249 1676 13252
rect 1664 13203 1676 13249
rect 1670 13200 1676 13203
rect 1728 13200 1734 13252
rect 2792 13181 2820 13348
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 3789 13311 3847 13317
rect 2924 13280 3372 13308
rect 2924 13268 2930 13280
rect 3344 13252 3372 13280
rect 3789 13277 3801 13311
rect 3835 13308 3847 13311
rect 3878 13308 3884 13320
rect 3835 13280 3884 13308
rect 3835 13277 3847 13280
rect 3789 13271 3847 13277
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4522 13308 4528 13320
rect 4111 13280 4528 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 3145 13243 3203 13249
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 3234 13240 3240 13252
rect 3191 13212 3240 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 3326 13200 3332 13252
rect 3384 13200 3390 13252
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 4080 13240 4108 13271
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 3752 13212 4108 13240
rect 3752 13200 3758 13212
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 2866 13172 2872 13184
rect 2823 13144 2872 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3881 13175 3939 13181
rect 3881 13172 3893 13175
rect 3016 13144 3893 13172
rect 3016 13132 3022 13144
rect 3881 13141 3893 13144
rect 3927 13141 3939 13175
rect 4632 13172 4660 13416
rect 4893 13413 4905 13447
rect 4939 13444 4951 13447
rect 5460 13444 5488 13472
rect 7852 13444 7880 13472
rect 4939 13416 5488 13444
rect 6564 13416 7880 13444
rect 4939 13413 4951 13416
rect 4893 13407 4951 13413
rect 4982 13336 4988 13388
rect 5040 13336 5046 13388
rect 6178 13336 6184 13388
rect 6236 13336 6242 13388
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5000 13308 5028 13336
rect 4939 13280 5028 13308
rect 5353 13321 5411 13327
rect 5353 13287 5365 13321
rect 5399 13287 5411 13321
rect 5353 13281 5411 13287
rect 6196 13308 6224 13336
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5368 13252 5396 13281
rect 6196 13280 6285 13308
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6564 13317 6592 13416
rect 8754 13336 8760 13388
rect 8812 13336 8818 13388
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 9548 13348 12112 13376
rect 9548 13336 9554 13348
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6420 13280 6561 13308
rect 6420 13268 6426 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 9766 13308 9772 13320
rect 9631 13280 9772 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 11330 13308 11336 13320
rect 9824 13280 11336 13308
rect 9824 13268 9830 13280
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11790 13268 11796 13320
rect 11848 13268 11854 13320
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12084 13317 12112 13348
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 13814 13308 13820 13320
rect 12115 13280 13820 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 5350 13200 5356 13252
rect 5408 13200 5414 13252
rect 8512 13243 8570 13249
rect 8512 13209 8524 13243
rect 8558 13240 8570 13243
rect 9398 13240 9404 13252
rect 8558 13212 9404 13240
rect 8558 13209 8570 13212
rect 8512 13203 8570 13209
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 5166 13172 5172 13184
rect 4632 13144 5172 13172
rect 3881 13135 3939 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5258 13132 5264 13184
rect 5316 13172 5322 13184
rect 5442 13172 5448 13184
rect 5316 13144 5448 13172
rect 5316 13132 5322 13144
rect 5442 13132 5448 13144
rect 5500 13172 5506 13184
rect 6365 13175 6423 13181
rect 6365 13172 6377 13175
rect 5500 13144 6377 13172
rect 5500 13132 5506 13144
rect 6365 13141 6377 13144
rect 6411 13141 6423 13175
rect 6365 13135 6423 13141
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 7466 13172 7472 13184
rect 7423 13144 7472 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 9214 13132 9220 13184
rect 9272 13132 9278 13184
rect 1104 13082 14536 13104
rect 1104 13030 4918 13082
rect 4970 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 5238 13082
rect 5290 13030 10918 13082
rect 10970 13030 10982 13082
rect 11034 13030 11046 13082
rect 11098 13030 11110 13082
rect 11162 13030 11174 13082
rect 11226 13030 11238 13082
rect 11290 13030 14536 13082
rect 1104 13008 14536 13030
rect 1670 12928 1676 12980
rect 1728 12928 1734 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5350 12968 5356 12980
rect 5123 12940 5356 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6236 12940 6377 12968
rect 6236 12928 6242 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 9490 12968 9496 12980
rect 6365 12931 6423 12937
rect 8956 12940 9496 12968
rect 4890 12860 4896 12912
rect 4948 12860 4954 12912
rect 6533 12903 6591 12909
rect 6533 12869 6545 12903
rect 6579 12900 6591 12903
rect 6579 12872 6684 12900
rect 6579 12869 6591 12872
rect 6533 12863 6591 12869
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 1857 12835 1915 12841
rect 1857 12832 1869 12835
rect 1728 12804 1869 12832
rect 1728 12792 1734 12804
rect 1857 12801 1869 12804
rect 1903 12801 1915 12835
rect 6656 12832 6684 12872
rect 6730 12860 6736 12912
rect 6788 12860 6794 12912
rect 8846 12832 8852 12844
rect 6656 12804 8852 12832
rect 1857 12795 1915 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 8956 12841 8984 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9732 12940 11652 12968
rect 9732 12928 9738 12940
rect 9861 12903 9919 12909
rect 9861 12900 9873 12903
rect 9416 12872 9873 12900
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9416 12841 9444 12872
rect 9861 12869 9873 12872
rect 9907 12869 9919 12903
rect 9861 12863 9919 12869
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 9180 12804 9413 12832
rect 9180 12792 9186 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 9784 12764 9812 12792
rect 9079 12736 9812 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 4522 12656 4528 12708
rect 4580 12656 4586 12708
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5684 12668 6592 12696
rect 5684 12656 5690 12668
rect 4614 12588 4620 12640
rect 4672 12628 4678 12640
rect 6564 12637 6592 12668
rect 4893 12631 4951 12637
rect 4893 12628 4905 12631
rect 4672 12600 4905 12628
rect 4672 12588 4678 12600
rect 4893 12597 4905 12600
rect 4939 12597 4951 12631
rect 4893 12591 4951 12597
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 8754 12588 8760 12640
rect 8812 12588 8818 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9968 12628 9996 12940
rect 10060 12872 10364 12900
rect 10060 12640 10088 12872
rect 10336 12841 10364 12872
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 11422 12832 11428 12844
rect 10321 12795 10379 12801
rect 10428 12804 11428 12832
rect 10244 12764 10272 12795
rect 10428 12764 10456 12804
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 10244 12736 10456 12764
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10560 12736 11529 12764
rect 10560 12724 10566 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11624 12764 11652 12940
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12897 12971 12955 12977
rect 12897 12968 12909 12971
rect 12492 12940 12909 12968
rect 12492 12928 12498 12940
rect 12897 12937 12909 12940
rect 12943 12937 12955 12971
rect 12897 12931 12955 12937
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13814 12968 13820 12980
rect 13587 12940 13820 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 11992 12900 12020 12928
rect 11808 12872 12020 12900
rect 11808 12841 11836 12872
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 11974 12832 11980 12844
rect 11931 12804 11980 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12084 12764 12112 12795
rect 11624 12736 12112 12764
rect 11517 12727 11575 12733
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 11790 12696 11796 12708
rect 11747 12668 11796 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 11790 12656 11796 12668
rect 11848 12656 11854 12708
rect 12084 12640 12112 12736
rect 13078 12724 13084 12776
rect 13136 12724 13142 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 9355 12600 9996 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 10042 12588 10048 12640
rect 10100 12588 10106 12640
rect 11606 12588 11612 12640
rect 11664 12588 11670 12640
rect 12066 12588 12072 12640
rect 12124 12588 12130 12640
rect 1104 12538 14536 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13918 12538
rect 13970 12486 13982 12538
rect 14034 12486 14046 12538
rect 14098 12486 14110 12538
rect 14162 12486 14174 12538
rect 14226 12486 14238 12538
rect 14290 12486 14536 12538
rect 1104 12464 14536 12486
rect 1670 12384 1676 12436
rect 1728 12384 1734 12436
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3510 12424 3516 12436
rect 2924 12396 3516 12424
rect 2924 12384 2930 12396
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4172 12396 4261 12424
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2961 12359 3019 12365
rect 2961 12356 2973 12359
rect 1903 12328 2973 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2961 12325 2973 12328
rect 3007 12325 3019 12359
rect 2961 12319 3019 12325
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2372 12260 2421 12288
rect 2372 12248 2378 12260
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2409 12251 2467 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3050 12288 3056 12300
rect 2823 12260 3056 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3050 12248 3056 12260
rect 3108 12288 3114 12300
rect 3237 12291 3295 12297
rect 3237 12288 3249 12291
rect 3108 12260 3249 12288
rect 3108 12248 3114 12260
rect 3237 12257 3249 12260
rect 3283 12257 3295 12291
rect 3237 12251 3295 12257
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3375 12260 4108 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 2498 12180 2504 12232
rect 2556 12180 2562 12232
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3142 12220 3148 12232
rect 2915 12192 3148 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 2133 12155 2191 12161
rect 2133 12121 2145 12155
rect 2179 12152 2191 12155
rect 2225 12155 2283 12161
rect 2225 12152 2237 12155
rect 2179 12124 2237 12152
rect 2179 12121 2191 12124
rect 2133 12115 2191 12121
rect 2225 12121 2237 12124
rect 2271 12121 2283 12155
rect 2225 12115 2283 12121
rect 2700 12124 2820 12152
rect 2700 12093 2728 12124
rect 2685 12087 2743 12093
rect 2685 12053 2697 12087
rect 2731 12053 2743 12087
rect 2792 12084 2820 12124
rect 3344 12084 3372 12251
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3510 12220 3516 12232
rect 3467 12192 3516 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 4080 12096 4108 12260
rect 2792 12056 3372 12084
rect 2685 12047 2743 12053
rect 4062 12044 4068 12096
rect 4120 12044 4126 12096
rect 4172 12084 4200 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 4249 12387 4307 12393
rect 4356 12396 4813 12424
rect 4233 12155 4291 12161
rect 4233 12121 4245 12155
rect 4279 12152 4291 12155
rect 4356 12152 4384 12396
rect 4801 12393 4813 12396
rect 4847 12424 4859 12427
rect 7009 12427 7067 12433
rect 4847 12396 6224 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 4430 12316 4436 12368
rect 4488 12356 4494 12368
rect 4706 12356 4712 12368
rect 4488 12328 4712 12356
rect 4488 12316 4494 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 6196 12365 6224 12396
rect 7009 12393 7021 12427
rect 7055 12424 7067 12427
rect 7098 12424 7104 12436
rect 7055 12396 7104 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7800 12396 7849 12424
rect 7800 12384 7806 12396
rect 7837 12393 7849 12396
rect 7883 12424 7895 12427
rect 8389 12427 8447 12433
rect 8389 12424 8401 12427
rect 7883 12396 8401 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 8389 12393 8401 12396
rect 8435 12424 8447 12427
rect 9214 12424 9220 12436
rect 8435 12396 9220 12424
rect 8435 12393 8447 12396
rect 8389 12387 8447 12393
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10744 12396 10977 12424
rect 10744 12384 10750 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 11425 12427 11483 12433
rect 10965 12387 11023 12393
rect 11072 12396 11376 12424
rect 6181 12359 6239 12365
rect 6181 12325 6193 12359
rect 6227 12356 6239 12359
rect 7377 12359 7435 12365
rect 7377 12356 7389 12359
rect 6227 12328 7389 12356
rect 6227 12325 6239 12328
rect 6181 12319 6239 12325
rect 7377 12325 7389 12328
rect 7423 12325 7435 12359
rect 9953 12359 10011 12365
rect 7377 12319 7435 12325
rect 7760 12328 8248 12356
rect 6730 12288 6736 12300
rect 4448 12260 6736 12288
rect 4448 12161 4476 12260
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7760 12297 7788 12328
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 7892 12260 8156 12288
rect 7892 12248 7898 12260
rect 5000 12192 6776 12220
rect 5000 12161 5028 12192
rect 4279 12124 4384 12152
rect 4433 12155 4491 12161
rect 4279 12121 4291 12124
rect 4233 12115 4291 12121
rect 4433 12121 4445 12155
rect 4479 12121 4491 12155
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4433 12115 4491 12121
rect 4540 12124 4997 12152
rect 4540 12084 4568 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 4985 12115 5043 12121
rect 5552 12124 5917 12152
rect 5552 12096 5580 12124
rect 5905 12121 5917 12124
rect 5951 12152 5963 12155
rect 5951 12124 6132 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 4172 12056 4568 12084
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 4785 12087 4843 12093
rect 4785 12053 4797 12087
rect 4831 12084 4843 12087
rect 5534 12084 5540 12096
rect 4831 12056 5540 12084
rect 4831 12053 4843 12056
rect 4785 12047 4843 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5626 12044 5632 12096
rect 5684 12044 5690 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 5813 12087 5871 12093
rect 5813 12084 5825 12087
rect 5776 12056 5825 12084
rect 5776 12044 5782 12056
rect 5813 12053 5825 12056
rect 5859 12053 5871 12087
rect 5813 12047 5871 12053
rect 5994 12044 6000 12096
rect 6052 12044 6058 12096
rect 6104 12084 6132 12124
rect 6641 12087 6699 12093
rect 6641 12084 6653 12087
rect 6104 12056 6653 12084
rect 6641 12053 6653 12056
rect 6687 12053 6699 12087
rect 6748 12084 6776 12192
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 7021 12223 7079 12229
rect 7021 12189 7033 12223
rect 7067 12220 7079 12223
rect 7067 12192 7420 12220
rect 7067 12189 7079 12192
rect 7021 12183 7079 12189
rect 7392 12152 7420 12192
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 7524 12192 7573 12220
rect 7524 12180 7530 12192
rect 7561 12189 7573 12192
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 8128 12229 8156 12260
rect 8220 12229 8248 12328
rect 9953 12325 9965 12359
rect 9999 12356 10011 12359
rect 10042 12356 10048 12368
rect 9999 12328 10048 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 11072 12288 11100 12396
rect 10744 12260 11100 12288
rect 10744 12248 10750 12260
rect 8113 12223 8171 12229
rect 7708 12192 7972 12220
rect 7708 12180 7714 12192
rect 7668 12152 7696 12180
rect 7392 12124 7696 12152
rect 7834 12112 7840 12164
rect 7892 12112 7898 12164
rect 7944 12152 7972 12192
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 8570 12220 8576 12232
rect 8251 12192 8576 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 10226 12220 10232 12232
rect 8904 12192 10232 12220
rect 8904 12180 8910 12192
rect 10226 12180 10232 12192
rect 10284 12220 10290 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10284 12192 10333 12220
rect 10284 12180 10290 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10857 12229 10885 12260
rect 11348 12239 11376 12396
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 12158 12424 12164 12436
rect 11471 12396 12164 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13136 12396 13645 12424
rect 13136 12384 13142 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12437 12359 12495 12365
rect 11572 12328 12204 12356
rect 11572 12316 11578 12328
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 11664 12260 12020 12288
rect 11664 12248 11670 12260
rect 11333 12233 11391 12239
rect 10827 12223 10885 12229
rect 10468 12192 10513 12220
rect 10468 12180 10474 12192
rect 10827 12189 10839 12223
rect 10873 12189 10885 12223
rect 10827 12183 10885 12189
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 7944 12124 8401 12152
rect 8389 12121 8401 12124
rect 8435 12152 8447 12155
rect 9306 12152 9312 12164
rect 8435 12124 9312 12152
rect 8435 12121 8447 12124
rect 8389 12115 8447 12121
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 9582 12112 9588 12164
rect 9640 12112 9646 12164
rect 10597 12155 10655 12161
rect 10597 12121 10609 12155
rect 10643 12121 10655 12155
rect 10597 12115 10655 12121
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 6748 12056 7941 12084
rect 6641 12047 6699 12053
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8076 12056 8585 12084
rect 8076 12044 8082 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 10042 12044 10048 12096
rect 10100 12044 10106 12096
rect 10612 12084 10640 12115
rect 10686 12112 10692 12164
rect 10744 12152 10750 12164
rect 11072 12152 11100 12183
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 11333 12199 11345 12233
rect 11379 12199 11391 12233
rect 11333 12193 11391 12199
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 10744 12124 11100 12152
rect 11149 12155 11207 12161
rect 10744 12112 10750 12124
rect 11149 12121 11161 12155
rect 11195 12152 11207 12155
rect 11532 12152 11560 12183
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 11992 12229 12020 12260
rect 12176 12229 12204 12328
rect 12437 12325 12449 12359
rect 12483 12356 12495 12359
rect 12526 12356 12532 12368
rect 12483 12328 12532 12356
rect 12483 12325 12495 12328
rect 12437 12319 12495 12325
rect 12526 12316 12532 12328
rect 12584 12356 12590 12368
rect 13170 12356 13176 12368
rect 12584 12328 13176 12356
rect 12584 12316 12590 12328
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 13872 12260 13952 12288
rect 13872 12248 13878 12260
rect 13924 12229 13952 12260
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11756 12192 11805 12220
rect 11756 12180 11762 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12220 12219 12223
rect 13909 12223 13967 12229
rect 12207 12192 12261 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 13909 12189 13921 12223
rect 13955 12189 13967 12223
rect 13909 12183 13967 12189
rect 12084 12152 12112 12183
rect 11195 12124 12112 12152
rect 12176 12152 12204 12183
rect 13265 12155 13323 12161
rect 13265 12152 13277 12155
rect 12176 12124 13277 12152
rect 11195 12121 11207 12124
rect 11149 12115 11207 12121
rect 13265 12121 13277 12124
rect 13311 12121 13323 12155
rect 13265 12115 13323 12121
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 13817 12155 13875 12161
rect 13817 12152 13829 12155
rect 13504 12124 13829 12152
rect 13504 12112 13510 12124
rect 13817 12121 13829 12124
rect 13863 12121 13875 12155
rect 13817 12115 13875 12121
rect 11790 12084 11796 12096
rect 10612 12056 11796 12084
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 1104 11994 14536 12016
rect 1104 11942 4918 11994
rect 4970 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 5238 11994
rect 5290 11942 10918 11994
rect 10970 11942 10982 11994
rect 11034 11942 11046 11994
rect 11098 11942 11110 11994
rect 11162 11942 11174 11994
rect 11226 11942 11238 11994
rect 11290 11942 14536 11994
rect 1104 11920 14536 11942
rect 3326 11840 3332 11892
rect 3384 11880 3390 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 3384 11852 4537 11880
rect 3384 11840 3390 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 4525 11843 4583 11849
rect 4693 11883 4751 11889
rect 4693 11849 4705 11883
rect 4739 11880 4751 11883
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4739 11852 4997 11880
rect 4739 11849 4751 11852
rect 4693 11843 4751 11849
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 5153 11883 5211 11889
rect 5153 11849 5165 11883
rect 5199 11880 5211 11883
rect 5442 11880 5448 11892
rect 5199 11852 5448 11880
rect 5199 11849 5211 11852
rect 5153 11843 5211 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5613 11883 5671 11889
rect 5613 11849 5625 11883
rect 5659 11880 5671 11883
rect 5718 11880 5724 11892
rect 5659 11852 5724 11880
rect 5659 11849 5671 11852
rect 5613 11843 5671 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 7282 11880 7288 11892
rect 7156 11852 7288 11880
rect 7156 11840 7162 11852
rect 7282 11840 7288 11852
rect 7340 11880 7346 11892
rect 8018 11880 8024 11892
rect 7340 11852 8024 11880
rect 7340 11840 7346 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 11422 11880 11428 11892
rect 9640 11852 11428 11880
rect 9640 11840 9646 11852
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 12066 11880 12072 11892
rect 11900 11852 12072 11880
rect 4890 11772 4896 11824
rect 4948 11772 4954 11824
rect 5258 11772 5264 11824
rect 5316 11812 5322 11824
rect 5353 11815 5411 11821
rect 5353 11812 5365 11815
rect 5316 11784 5365 11812
rect 5316 11772 5322 11784
rect 5353 11781 5365 11784
rect 5399 11781 5411 11815
rect 5353 11775 5411 11781
rect 5810 11772 5816 11824
rect 5868 11772 5874 11824
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 11790 11812 11796 11824
rect 10827 11784 11796 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4430 11704 4436 11756
rect 4488 11704 4494 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 8536 11716 8585 11744
rect 8536 11704 8542 11716
rect 8573 11713 8585 11716
rect 8619 11744 8631 11747
rect 9122 11744 9128 11756
rect 8619 11716 9128 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 9416 11716 10701 11744
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 4448 11676 4476 11704
rect 9416 11676 9444 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11256 11716 11529 11744
rect 11256 11676 11284 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11900 11753 11928 11852
rect 12066 11840 12072 11852
rect 12124 11880 12130 11892
rect 12124 11852 12664 11880
rect 12124 11840 12130 11852
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 12250 11704 12256 11756
rect 12308 11704 12314 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 3835 11648 4476 11676
rect 8956 11648 9444 11676
rect 10428 11648 11284 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 5445 11611 5503 11617
rect 5445 11608 5457 11611
rect 4816 11580 5457 11608
rect 4816 11552 4844 11580
rect 5445 11577 5457 11580
rect 5491 11577 5503 11611
rect 5445 11571 5503 11577
rect 8956 11552 8984 11648
rect 10428 11552 10456 11648
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11388 11648 11713 11676
rect 11388 11636 11394 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 12452 11676 12480 11707
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12636 11744 12664 11852
rect 13446 11840 13452 11892
rect 13504 11840 13510 11892
rect 12986 11772 12992 11824
rect 13044 11812 13050 11824
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 13044 11784 13553 11812
rect 13044 11772 13050 11784
rect 13541 11781 13553 11784
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12636 11716 12817 11744
rect 12805 11713 12817 11716
rect 12851 11744 12863 11747
rect 13814 11744 13820 11756
rect 12851 11716 13820 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 11701 11639 11759 11645
rect 11900 11648 12480 11676
rect 12621 11679 12679 11685
rect 10502 11568 10508 11620
rect 10560 11568 10566 11620
rect 11900 11617 11928 11648
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12894 11676 12900 11688
rect 12621 11639 12679 11645
rect 12717 11648 12900 11676
rect 11885 11611 11943 11617
rect 11885 11577 11897 11611
rect 11931 11577 11943 11611
rect 11885 11571 11943 11577
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12636 11608 12664 11639
rect 12216 11580 12664 11608
rect 12216 11568 12222 11580
rect 4154 11500 4160 11552
rect 4212 11500 4218 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4614 11540 4620 11552
rect 4396 11512 4620 11540
rect 4396 11500 4402 11512
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 4798 11540 4804 11552
rect 4755 11512 4804 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5534 11540 5540 11552
rect 5215 11512 5540 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5902 11540 5908 11552
rect 5675 11512 5908 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 8938 11540 8944 11552
rect 8803 11512 8944 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 10410 11500 10416 11552
rect 10468 11500 10474 11552
rect 10520 11540 10548 11568
rect 12717 11540 12745 11648
rect 12894 11636 12900 11648
rect 12952 11676 12958 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12952 11648 13185 11676
rect 12952 11636 12958 11648
rect 13173 11645 13185 11648
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 12989 11611 13047 11617
rect 12989 11577 13001 11611
rect 13035 11608 13047 11611
rect 13265 11611 13323 11617
rect 13265 11608 13277 11611
rect 13035 11580 13277 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 13265 11577 13277 11580
rect 13311 11577 13323 11611
rect 13265 11571 13323 11577
rect 10520 11512 12745 11540
rect 13078 11500 13084 11552
rect 13136 11500 13142 11552
rect 1104 11450 14536 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13918 11450
rect 13970 11398 13982 11450
rect 14034 11398 14046 11450
rect 14098 11398 14110 11450
rect 14162 11398 14174 11450
rect 14226 11398 14238 11450
rect 14290 11398 14536 11450
rect 1104 11376 14536 11398
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3200 11308 3801 11336
rect 3200 11296 3206 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4154 11296 4160 11348
rect 4212 11296 4218 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 5868 11308 8309 11336
rect 5868 11296 5874 11308
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 8803 11308 9076 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 1949 11271 2007 11277
rect 1949 11237 1961 11271
rect 1995 11268 2007 11271
rect 2317 11271 2375 11277
rect 2317 11268 2329 11271
rect 1995 11240 2329 11268
rect 1995 11237 2007 11240
rect 1949 11231 2007 11237
rect 2317 11237 2329 11240
rect 2363 11237 2375 11271
rect 2317 11231 2375 11237
rect 1762 11160 1768 11212
rect 1820 11160 1826 11212
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2866 11200 2872 11212
rect 2547 11172 2872 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 2222 11024 2228 11076
rect 2280 11024 2286 11076
rect 2608 11064 2636 11095
rect 2682 11092 2688 11144
rect 2740 11092 2746 11144
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 2958 11132 2964 11144
rect 2823 11104 2964 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 2958 11092 2964 11104
rect 3016 11132 3022 11144
rect 3602 11132 3608 11144
rect 3016 11104 3608 11132
rect 3016 11092 3022 11104
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3844 11104 4077 11132
rect 3844 11092 3850 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4172 11132 4200 11296
rect 4890 11268 4896 11280
rect 4356 11240 4896 11268
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 4172 11104 4261 11132
rect 4065 11095 4123 11101
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 4356 11132 4384 11240
rect 4890 11228 4896 11240
rect 4948 11228 4954 11280
rect 6730 11268 6736 11280
rect 5276 11240 6736 11268
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4798 11200 4804 11212
rect 4479 11172 4804 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 4525 11135 4583 11141
rect 4356 11104 4476 11132
rect 4249 11095 4307 11101
rect 4338 11064 4344 11076
rect 2608 11036 4344 11064
rect 2700 11008 2728 11036
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 2682 10956 2688 11008
rect 2740 10956 2746 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4157 10999 4215 11005
rect 4157 10996 4169 10999
rect 4028 10968 4169 10996
rect 4028 10956 4034 10968
rect 4157 10965 4169 10968
rect 4203 10996 4215 10999
rect 4448 10996 4476 11104
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4890 11132 4896 11144
rect 4571 11104 4896 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5276 11141 5304 11240
rect 6730 11228 6736 11240
rect 6788 11268 6794 11280
rect 7469 11271 7527 11277
rect 7469 11268 7481 11271
rect 6788 11240 7481 11268
rect 6788 11228 6794 11240
rect 7469 11237 7481 11240
rect 7515 11237 7527 11271
rect 7469 11231 7527 11237
rect 7558 11228 7564 11280
rect 7616 11228 7622 11280
rect 7742 11228 7748 11280
rect 7800 11228 7806 11280
rect 9048 11277 9076 11308
rect 9398 11296 9404 11348
rect 9456 11296 9462 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 12986 11336 12992 11348
rect 10284 11308 12992 11336
rect 10284 11296 10290 11308
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 9214 11268 9220 11280
rect 9079 11240 9220 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 10134 11268 10140 11280
rect 9916 11240 10140 11268
rect 9916 11228 9922 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 5736 11172 6285 11200
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 5000 11064 5028 11095
rect 4856 11036 5028 11064
rect 5092 11064 5120 11095
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 5736 11141 5764 11172
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 6914 11200 6920 11212
rect 6273 11163 6331 11169
rect 6472 11172 6684 11200
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 5500 11104 5733 11132
rect 5500 11092 5506 11104
rect 5721 11101 5733 11104
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 5828 11064 5856 11095
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 5994 11092 6000 11144
rect 6052 11092 6058 11144
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6472 11132 6500 11172
rect 6656 11144 6684 11172
rect 6748 11172 6920 11200
rect 6227 11104 6500 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 6638 11092 6644 11144
rect 6696 11092 6702 11144
rect 6748 11141 6776 11172
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7576 11200 7604 11228
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 6972 11172 7144 11200
rect 7576 11172 7849 11200
rect 6972 11160 6978 11172
rect 7116 11144 7144 11172
rect 7837 11169 7849 11172
rect 7883 11200 7895 11203
rect 7883 11172 8156 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6822 11092 6828 11144
rect 6880 11092 6886 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 6914 11064 6920 11076
rect 5092 11036 5580 11064
rect 5828 11036 6920 11064
rect 4856 11024 4862 11036
rect 4203 10968 4476 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 4614 10956 4620 11008
rect 4672 10956 4678 11008
rect 5000 10996 5028 11036
rect 5258 10996 5264 11008
rect 5000 10968 5264 10996
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 5552 10996 5580 11036
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 7024 11064 7052 11095
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7926 11132 7932 11144
rect 7156 11104 7932 11132
rect 7156 11092 7162 11104
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 7650 11064 7656 11076
rect 7024 11036 7656 11064
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 8128 11064 8156 11172
rect 8220 11172 8616 11200
rect 8220 11141 8248 11172
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8478 11132 8484 11144
rect 8205 11095 8263 11101
rect 8404 11104 8484 11132
rect 8404 11064 8432 11104
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8588 11132 8616 11172
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9490 11200 9496 11212
rect 8996 11172 9496 11200
rect 8996 11160 9002 11172
rect 9490 11160 9496 11172
rect 9548 11200 9554 11212
rect 11330 11200 11336 11212
rect 9548 11172 9720 11200
rect 9548 11160 9554 11172
rect 8588 11104 8800 11132
rect 8772 11076 8800 11104
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9692 11141 9720 11172
rect 9784 11172 11336 11200
rect 9784 11144 9812 11172
rect 11330 11160 11336 11172
rect 11388 11200 11394 11212
rect 11698 11200 11704 11212
rect 11388 11172 11704 11200
rect 11388 11160 11394 11172
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 9180 11104 9229 11132
rect 9180 11092 9186 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10134 11132 10140 11144
rect 10091 11104 10140 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 10134 11092 10140 11104
rect 10192 11132 10198 11144
rect 10192 11104 10916 11132
rect 10192 11092 10198 11104
rect 8128 11036 8432 11064
rect 8754 11024 8760 11076
rect 8812 11024 8818 11076
rect 10778 11024 10784 11076
rect 10836 11024 10842 11076
rect 10888 11064 10916 11104
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11790 11132 11796 11144
rect 11112 11104 11796 11132
rect 11112 11092 11118 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 10888 11036 11928 11064
rect 11900 11008 11928 11036
rect 5718 10996 5724 11008
rect 5552 10968 5724 10996
rect 5718 10956 5724 10968
rect 5776 10996 5782 11008
rect 6454 10996 6460 11008
rect 5776 10968 6460 10996
rect 5776 10956 5782 10968
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 8113 10999 8171 11005
rect 8113 10996 8125 10999
rect 6788 10968 8125 10996
rect 6788 10956 6794 10968
rect 8113 10965 8125 10968
rect 8159 10965 8171 10999
rect 8113 10959 8171 10965
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 10686 10996 10692 11008
rect 9088 10968 10692 10996
rect 9088 10956 9094 10968
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11882 10956 11888 11008
rect 11940 10956 11946 11008
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 12526 10996 12532 11008
rect 12299 10968 12532 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12526 10956 12532 10968
rect 12584 10996 12590 11008
rect 12710 10996 12716 11008
rect 12584 10968 12716 10996
rect 12584 10956 12590 10968
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 1104 10906 14536 10928
rect 1104 10854 4918 10906
rect 4970 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 5238 10906
rect 5290 10854 10918 10906
rect 10970 10854 10982 10906
rect 11034 10854 11046 10906
rect 11098 10854 11110 10906
rect 11162 10854 11174 10906
rect 11226 10854 11238 10906
rect 11290 10854 14536 10906
rect 1104 10832 14536 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2222 10792 2228 10804
rect 2179 10764 2228 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 2222 10752 2228 10764
rect 2280 10752 2286 10804
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10761 2651 10795
rect 2593 10755 2651 10761
rect 2608 10724 2636 10755
rect 2682 10752 2688 10804
rect 2740 10752 2746 10804
rect 2774 10752 2780 10804
rect 2832 10752 2838 10804
rect 3878 10752 3884 10804
rect 3936 10752 3942 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4614 10792 4620 10804
rect 4019 10764 4620 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5442 10792 5448 10804
rect 5307 10764 5448 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8662 10792 8668 10804
rect 7984 10764 8668 10792
rect 7984 10752 7990 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 9030 10752 9036 10804
rect 9088 10752 9094 10804
rect 9585 10795 9643 10801
rect 9585 10761 9597 10795
rect 9631 10792 9643 10795
rect 9858 10792 9864 10804
rect 9631 10764 9864 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10792 10471 10795
rect 10686 10792 10692 10804
rect 10459 10764 10692 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 11146 10792 11152 10804
rect 11204 10801 11210 10804
rect 11204 10795 11223 10801
rect 10928 10764 11152 10792
rect 10928 10752 10934 10764
rect 11146 10752 11152 10764
rect 11211 10761 11223 10795
rect 11204 10755 11223 10761
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11606 10792 11612 10804
rect 11379 10764 11612 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11204 10752 11210 10755
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13872 10764 13921 10792
rect 13872 10752 13878 10764
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 13909 10755 13967 10761
rect 2792 10724 2820 10752
rect 2608 10696 2820 10724
rect 3896 10724 3924 10752
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 3896 10696 5089 10724
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2590 10656 2596 10668
rect 2372 10628 2596 10656
rect 2372 10616 2378 10628
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2498 10588 2504 10600
rect 2455 10560 2504 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2700 10588 2728 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5353 10727 5411 10733
rect 5353 10693 5365 10727
rect 5399 10724 5411 10727
rect 5626 10724 5632 10736
rect 5399 10696 5632 10724
rect 5399 10693 5411 10696
rect 5353 10687 5411 10693
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 9401 10727 9459 10733
rect 5960 10696 6776 10724
rect 5960 10684 5966 10696
rect 6748 10668 6776 10696
rect 6932 10696 7328 10724
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2866 10656 2872 10668
rect 2823 10628 2872 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2866 10616 2872 10628
rect 2924 10656 2930 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 2924 10628 3525 10656
rect 2924 10616 2930 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 3786 10616 3792 10668
rect 3844 10616 3850 10668
rect 3878 10616 3884 10668
rect 3936 10616 3942 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4798 10656 4804 10668
rect 4203 10628 4804 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 4856 10628 5457 10656
rect 4856 10616 4862 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6546 10656 6552 10668
rect 6052 10628 6552 10656
rect 6052 10616 6058 10628
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 3050 10588 3056 10600
rect 2700 10560 3056 10588
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3804 10452 3832 10616
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4338 10588 4344 10600
rect 4295 10560 4344 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 6656 10588 6684 10619
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 6932 10665 6960 10696
rect 7300 10668 7328 10696
rect 9401 10693 9413 10727
rect 9447 10724 9459 10727
rect 9447 10696 10364 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7098 10656 7104 10668
rect 7055 10628 7104 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8628 10628 8677 10656
rect 8628 10616 8634 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9355 10628 9444 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 7190 10588 7196 10600
rect 6656 10560 7196 10588
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 8496 10588 8524 10616
rect 9416 10600 9444 10628
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9692 10628 9781 10656
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8496 10560 8769 10588
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 5500 10492 5641 10520
rect 5500 10480 5506 10492
rect 5629 10489 5641 10492
rect 5675 10520 5687 10523
rect 5675 10492 7052 10520
rect 5675 10489 5687 10492
rect 5629 10483 5687 10489
rect 7024 10464 7052 10492
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 9692 10520 9720 10628
rect 9769 10625 9781 10628
rect 9815 10656 9827 10659
rect 10134 10656 10140 10668
rect 9815 10628 10140 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10336 10665 10364 10696
rect 10962 10684 10968 10736
rect 11020 10684 11026 10736
rect 11514 10724 11520 10736
rect 11072 10696 11520 10724
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 11072 10656 11100 10696
rect 11514 10684 11520 10696
rect 11572 10684 11578 10736
rect 11624 10724 11652 10752
rect 12796 10727 12854 10733
rect 11624 10696 11928 10724
rect 10643 10628 11100 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10244 10588 10272 10619
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11698 10656 11704 10668
rect 11480 10628 11704 10656
rect 11480 10616 11486 10628
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11900 10665 11928 10696
rect 12796 10693 12808 10727
rect 12842 10724 12854 10727
rect 13078 10724 13084 10736
rect 12842 10696 13084 10724
rect 12842 10693 12854 10696
rect 12796 10687 12854 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12250 10656 12256 10668
rect 12023 10628 12256 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 13722 10656 13728 10668
rect 12308 10628 13728 10656
rect 12308 10616 12314 10628
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 9999 10560 10088 10588
rect 10244 10560 11529 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 9180 10492 9720 10520
rect 9180 10480 9186 10492
rect 4246 10452 4252 10464
rect 3804 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 7006 10412 7012 10464
rect 7064 10412 7070 10464
rect 8846 10412 8852 10464
rect 8904 10412 8910 10464
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10060 10452 10088 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11808 10588 11836 10616
rect 11808 10560 11928 10588
rect 11517 10551 11575 10557
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 10888 10492 11805 10520
rect 10888 10464 10916 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 11793 10483 11851 10489
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 10060 10424 10609 10452
rect 10597 10421 10609 10424
rect 10643 10421 10655 10455
rect 10597 10415 10655 10421
rect 10870 10412 10876 10464
rect 10928 10412 10934 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10452 11207 10455
rect 11900 10452 11928 10560
rect 12526 10548 12532 10600
rect 12584 10548 12590 10600
rect 11195 10424 11928 10452
rect 12544 10452 12572 10548
rect 12802 10452 12808 10464
rect 12544 10424 12808 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 1104 10362 14536 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13918 10362
rect 13970 10310 13982 10362
rect 14034 10310 14046 10362
rect 14098 10310 14110 10362
rect 14162 10310 14174 10362
rect 14226 10310 14238 10362
rect 14290 10310 14536 10362
rect 1104 10288 14536 10310
rect 4433 10251 4491 10257
rect 4433 10217 4445 10251
rect 4479 10248 4491 10251
rect 4798 10248 4804 10260
rect 4479 10220 4804 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6604 10220 6837 10248
rect 6604 10208 6610 10220
rect 6825 10217 6837 10220
rect 6871 10248 6883 10251
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 6871 10220 7573 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 7561 10217 7573 10220
rect 7607 10248 7619 10251
rect 9214 10248 9220 10260
rect 7607 10220 9220 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 10870 10208 10876 10260
rect 10928 10208 10934 10260
rect 13722 10208 13728 10260
rect 13780 10208 13786 10260
rect 2777 10183 2835 10189
rect 2777 10149 2789 10183
rect 2823 10180 2835 10183
rect 2958 10180 2964 10192
rect 2823 10152 2964 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 2958 10140 2964 10152
rect 3016 10180 3022 10192
rect 3016 10152 6500 10180
rect 3016 10140 3022 10152
rect 4617 10115 4675 10121
rect 4617 10112 4629 10115
rect 3344 10084 4629 10112
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 1486 10044 1492 10056
rect 1443 10016 1492 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1486 10004 1492 10016
rect 1544 10044 1550 10056
rect 3344 10044 3372 10084
rect 4617 10081 4629 10084
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 6472 10056 6500 10152
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7745 10183 7803 10189
rect 7745 10180 7757 10183
rect 7064 10152 7757 10180
rect 7064 10140 7070 10152
rect 7745 10149 7757 10152
rect 7791 10149 7803 10183
rect 7745 10143 7803 10149
rect 8570 10140 8576 10192
rect 8628 10180 8634 10192
rect 11146 10180 11152 10192
rect 8628 10152 11152 10180
rect 8628 10140 8634 10152
rect 11146 10140 11152 10152
rect 11204 10140 11210 10192
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6696 10084 6745 10112
rect 6696 10072 6702 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 1544 10016 3372 10044
rect 1544 10004 1550 10016
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4396 10016 4537 10044
rect 4396 10004 4402 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6748 10044 6776 10075
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7469 10115 7527 10121
rect 6972 10084 7328 10112
rect 6972 10072 6978 10084
rect 6748 10016 7144 10044
rect 1664 9979 1722 9985
rect 1664 9945 1676 9979
rect 1710 9976 1722 9979
rect 1762 9976 1768 9988
rect 1710 9948 1768 9976
rect 1710 9945 1722 9948
rect 1664 9939 1722 9945
rect 1762 9936 1768 9948
rect 1820 9936 1826 9988
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 4157 9979 4215 9985
rect 4157 9976 4169 9979
rect 3936 9948 4169 9976
rect 3936 9936 3942 9948
rect 4157 9945 4169 9948
rect 4203 9976 4215 9979
rect 6365 9979 6423 9985
rect 4203 9948 4384 9976
rect 4203 9945 4215 9948
rect 4157 9939 4215 9945
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3384 9880 3801 9908
rect 3384 9868 3390 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 4246 9868 4252 9920
rect 4304 9868 4310 9920
rect 4356 9908 4384 9948
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 7116 9976 7144 10016
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7300 10053 7328 10084
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7834 10112 7840 10124
rect 7515 10084 7840 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8938 10112 8944 10124
rect 8036 10084 8944 10112
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 8036 10044 8064 10084
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 7607 10016 8064 10044
rect 8128 10016 8217 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 7576 9976 7604 10007
rect 8128 9988 8156 10016
rect 8205 10013 8217 10016
rect 8251 10044 8263 10047
rect 8570 10044 8576 10056
rect 8251 10016 8576 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8956 10044 8984 10072
rect 8956 10038 10829 10044
rect 10870 10038 10876 10056
rect 8956 10016 10876 10038
rect 10801 10010 10876 10016
rect 10870 10004 10876 10010
rect 10928 10004 10934 10056
rect 11164 10053 11192 10140
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11388 10084 12296 10112
rect 11388 10072 11394 10084
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10044 11207 10047
rect 11195 10016 12112 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 6411 9948 6868 9976
rect 7116 9948 7604 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 6840 9920 6868 9948
rect 8110 9936 8116 9988
rect 8168 9936 8174 9988
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9976 8355 9979
rect 8386 9976 8392 9988
rect 8343 9948 8392 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 8386 9936 8392 9948
rect 8444 9976 8450 9988
rect 12084 9976 12112 10016
rect 12158 10004 12164 10056
rect 12216 10004 12222 10056
rect 12268 10044 12296 10084
rect 12342 10044 12348 10056
rect 12268 10016 12348 10044
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 12434 9976 12440 9988
rect 8444 9948 11560 9976
rect 12084 9948 12440 9976
rect 8444 9936 8450 9948
rect 11532 9920 11560 9948
rect 12434 9936 12440 9948
rect 12492 9976 12498 9988
rect 12805 9979 12863 9985
rect 12805 9976 12817 9979
rect 12492 9948 12817 9976
rect 12492 9936 12498 9948
rect 12805 9945 12817 9948
rect 12851 9945 12863 9979
rect 12805 9939 12863 9945
rect 13170 9936 13176 9988
rect 13228 9936 13234 9988
rect 13354 9936 13360 9988
rect 13412 9936 13418 9988
rect 13541 9979 13599 9985
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13630 9976 13636 9988
rect 13587 9948 13636 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 4356 9880 6469 9908
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 6822 9868 6828 9920
rect 6880 9868 6886 9920
rect 7101 9911 7159 9917
rect 7101 9877 7113 9911
rect 7147 9908 7159 9911
rect 8202 9908 8208 9920
rect 7147 9880 8208 9908
rect 7147 9877 7159 9880
rect 7101 9871 7159 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 11054 9908 11060 9920
rect 9548 9880 11060 9908
rect 9548 9868 9554 9880
rect 11054 9868 11060 9880
rect 11112 9908 11118 9920
rect 11422 9908 11428 9920
rect 11112 9880 11428 9908
rect 11112 9868 11118 9880
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11514 9868 11520 9920
rect 11572 9868 11578 9920
rect 12250 9868 12256 9920
rect 12308 9868 12314 9920
rect 1104 9818 14536 9840
rect 1104 9766 4918 9818
rect 4970 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 5238 9818
rect 5290 9766 10918 9818
rect 10970 9766 10982 9818
rect 11034 9766 11046 9818
rect 11098 9766 11110 9818
rect 11162 9766 11174 9818
rect 11226 9766 11238 9818
rect 11290 9766 14536 9818
rect 1104 9744 14536 9766
rect 1762 9664 1768 9716
rect 1820 9664 1826 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4304 9676 4997 9704
rect 4304 9664 4310 9676
rect 4985 9673 4997 9676
rect 5031 9704 5043 9707
rect 5442 9704 5448 9716
rect 5031 9676 5448 9704
rect 5031 9673 5043 9676
rect 4985 9667 5043 9673
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5592 9676 7328 9704
rect 5592 9664 5598 9676
rect 1854 9596 1860 9648
rect 1912 9596 1918 9648
rect 4614 9636 4620 9648
rect 4080 9608 4620 9636
rect 1872 9568 1900 9596
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1872 9540 1961 9568
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 3142 9528 3148 9580
rect 3200 9568 3206 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3200 9540 3985 9568
rect 3200 9528 3206 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 3068 9500 3096 9528
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 3068 9472 3249 9500
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 3326 9460 3332 9512
rect 3384 9460 3390 9512
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3878 9500 3884 9512
rect 3467 9472 3884 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3878 9460 3884 9472
rect 3936 9500 3942 9512
rect 4080 9500 4108 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4798 9596 4804 9648
rect 4856 9636 4862 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4856 9608 4905 9636
rect 4856 9596 4862 9608
rect 4893 9605 4905 9608
rect 4939 9636 4951 9639
rect 5353 9639 5411 9645
rect 5353 9636 5365 9639
rect 4939 9608 5365 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 5353 9605 5365 9608
rect 5399 9605 5411 9639
rect 5353 9599 5411 9605
rect 5920 9608 6592 9636
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4338 9568 4344 9580
rect 4203 9540 4344 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 5626 9568 5632 9580
rect 4479 9540 5632 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5718 9528 5724 9580
rect 5776 9577 5782 9580
rect 5776 9571 5808 9577
rect 5796 9568 5808 9571
rect 5920 9568 5948 9608
rect 5796 9540 5948 9568
rect 5796 9537 5808 9540
rect 5776 9531 5808 9537
rect 5776 9528 5782 9531
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6089 9571 6147 9577
rect 6089 9568 6101 9571
rect 6052 9540 6101 9568
rect 6052 9528 6058 9540
rect 6089 9537 6101 9540
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 3936 9472 4108 9500
rect 3936 9460 3942 9472
rect 4614 9460 4620 9512
rect 4672 9460 4678 9512
rect 5102 9503 5160 9509
rect 5102 9469 5114 9503
rect 5148 9500 5160 9503
rect 6564 9500 6592 9608
rect 6914 9596 6920 9648
rect 6972 9596 6978 9648
rect 7300 9636 7328 9676
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 7834 9704 7840 9716
rect 7432 9676 7840 9704
rect 7432 9664 7438 9676
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 10778 9664 10784 9716
rect 10836 9664 10842 9716
rect 11793 9707 11851 9713
rect 11793 9673 11805 9707
rect 11839 9704 11851 9707
rect 12158 9704 12164 9716
rect 11839 9676 12164 9704
rect 11839 9673 11851 9676
rect 11793 9667 11851 9673
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12250 9664 12256 9716
rect 12308 9664 12314 9716
rect 12342 9664 12348 9716
rect 12400 9664 12406 9716
rect 8110 9636 8116 9648
rect 7300 9608 8116 9636
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 7190 9568 7196 9580
rect 6779 9540 7196 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7484 9577 7512 9608
rect 8110 9596 8116 9608
rect 8168 9596 8174 9648
rect 9398 9596 9404 9648
rect 9456 9636 9462 9648
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 9456 9608 10425 9636
rect 9456 9596 9462 9608
rect 10413 9605 10425 9608
rect 10459 9605 10471 9639
rect 10796 9636 10824 9664
rect 10796 9608 11376 9636
rect 10413 9599 10471 9605
rect 11348 9580 11376 9608
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 8803 9540 9321 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9309 9537 9321 9540
rect 9355 9568 9367 9571
rect 10597 9571 10655 9577
rect 9355 9540 10272 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 7300 9500 7328 9531
rect 7852 9500 7880 9531
rect 8846 9500 8852 9512
rect 5148 9472 5672 9500
rect 5148 9469 5160 9472
rect 5102 9463 5160 9469
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2866 9432 2872 9444
rect 2556 9404 2872 9432
rect 2556 9392 2562 9404
rect 2866 9392 2872 9404
rect 2924 9432 2930 9444
rect 4062 9432 4068 9444
rect 2924 9404 4068 9432
rect 2924 9392 2930 9404
rect 4062 9392 4068 9404
rect 4120 9432 4126 9444
rect 4249 9435 4307 9441
rect 4249 9432 4261 9435
rect 4120 9404 4261 9432
rect 4120 9392 4126 9404
rect 4249 9401 4261 9404
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 4341 9435 4399 9441
rect 4341 9401 4353 9435
rect 4387 9432 4399 9435
rect 4798 9432 4804 9444
rect 4387 9404 4804 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4798 9392 4804 9404
rect 4856 9392 4862 9444
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5350 9432 5356 9444
rect 5307 9404 5356 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 5644 9432 5672 9472
rect 5828 9472 6500 9500
rect 6564 9472 8852 9500
rect 5828 9432 5856 9472
rect 5644 9404 5856 9432
rect 5951 9435 6009 9441
rect 5951 9401 5963 9435
rect 5997 9432 6009 9435
rect 5997 9404 6224 9432
rect 5997 9401 6009 9404
rect 5951 9395 6009 9401
rect 6196 9376 6224 9404
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 6086 9364 6092 9376
rect 5859 9336 6092 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6178 9324 6184 9376
rect 6236 9324 6242 9376
rect 6472 9373 6500 9472
rect 8846 9460 8852 9472
rect 8904 9500 8910 9512
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 8904 9472 9045 9500
rect 8904 9460 8910 9472
rect 9033 9469 9045 9472
rect 9079 9500 9091 9503
rect 9490 9500 9496 9512
rect 9079 9472 9496 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 10244 9432 10272 9540
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10686 9568 10692 9580
rect 10643 9540 10692 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10796 9432 10824 9531
rect 11330 9528 11336 9580
rect 11388 9528 11394 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12268 9577 12296 9664
rect 12360 9577 12388 9664
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 11940 9540 12081 9568
rect 11940 9528 11946 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 12434 9528 12440 9580
rect 12492 9528 12498 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 13061 9571 13119 9577
rect 13061 9568 13073 9571
rect 12912 9540 13073 9568
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12526 9500 12532 9512
rect 11839 9472 12532 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12912 9500 12940 9540
rect 13061 9537 13073 9540
rect 13107 9537 13119 9571
rect 13061 9531 13119 9537
rect 12728 9472 12940 9500
rect 12728 9441 12756 9472
rect 12713 9435 12771 9441
rect 10244 9404 12434 9432
rect 6457 9367 6515 9373
rect 6457 9333 6469 9367
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 6604 9336 6653 9364
rect 6604 9324 6610 9336
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8386 9364 8392 9376
rect 8343 9336 8392 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 8754 9364 8760 9376
rect 8536 9336 8760 9364
rect 8536 9324 8542 9336
rect 8754 9324 8760 9336
rect 8812 9364 8818 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8812 9336 8953 9364
rect 8812 9324 8818 9336
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 8941 9327 8999 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 10008 9336 11621 9364
rect 10008 9324 10014 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 12406 9364 12434 9404
rect 12713 9401 12725 9435
rect 12759 9401 12771 9435
rect 12713 9395 12771 9401
rect 13170 9364 13176 9376
rect 12406 9336 13176 9364
rect 11609 9327 11667 9333
rect 13170 9324 13176 9336
rect 13228 9364 13234 9376
rect 14185 9367 14243 9373
rect 14185 9364 14197 9367
rect 13228 9336 14197 9364
rect 13228 9324 13234 9336
rect 14185 9333 14197 9336
rect 14231 9333 14243 9367
rect 14185 9327 14243 9333
rect 1104 9274 14536 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13918 9274
rect 13970 9222 13982 9274
rect 14034 9222 14046 9274
rect 14098 9222 14110 9274
rect 14162 9222 14174 9274
rect 14226 9222 14238 9274
rect 14290 9222 14536 9274
rect 1104 9200 14536 9222
rect 2958 9160 2964 9172
rect 2746 9132 2964 9160
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2746 9092 2774 9132
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 3142 9120 3148 9172
rect 3200 9120 3206 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 5442 9160 5448 9172
rect 4396 9132 5448 9160
rect 4396 9120 4402 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 6914 9160 6920 9172
rect 6135 9132 6920 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 9122 9160 9128 9172
rect 8260 9132 9128 9160
rect 8260 9120 8266 9132
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 12802 9160 12808 9172
rect 9876 9132 12808 9160
rect 2455 9064 2774 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2866 8984 2872 9036
rect 2924 8984 2930 9036
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 3160 9024 3188 9120
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 8757 9095 8815 9101
rect 7248 9064 8524 9092
rect 7248 9052 7254 9064
rect 3237 9027 3295 9033
rect 3237 9024 3249 9027
rect 3160 8996 3249 9024
rect 3237 8993 3249 8996
rect 3283 8993 3295 9027
rect 3237 8987 3295 8993
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 4614 9024 4620 9036
rect 3881 8987 3939 8993
rect 4172 8996 4620 9024
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2777 8959 2835 8965
rect 2777 8956 2789 8959
rect 2740 8928 2789 8956
rect 2740 8916 2746 8928
rect 2777 8925 2789 8928
rect 2823 8956 2835 8959
rect 2958 8956 2964 8968
rect 2823 8928 2964 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3068 8956 3096 8984
rect 3145 8959 3203 8965
rect 3145 8956 3157 8959
rect 3068 8928 3157 8956
rect 3145 8925 3157 8928
rect 3191 8956 3203 8959
rect 3896 8956 3924 8987
rect 4172 8965 4200 8996
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 4672 8996 6469 9024
rect 4672 8984 4678 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6840 8996 7052 9024
rect 3191 8928 3924 8956
rect 4157 8959 4215 8965
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6420 8928 6653 8956
rect 6420 8916 6426 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 2041 8891 2099 8897
rect 2041 8857 2053 8891
rect 2087 8888 2099 8891
rect 2593 8891 2651 8897
rect 2593 8888 2605 8891
rect 2087 8860 2605 8888
rect 2087 8857 2099 8860
rect 2041 8851 2099 8857
rect 2593 8857 2605 8860
rect 2639 8857 2651 8891
rect 2593 8851 2651 8857
rect 5721 8891 5779 8897
rect 5721 8857 5733 8891
rect 5767 8888 5779 8891
rect 5810 8888 5816 8900
rect 5767 8860 5816 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 5905 8891 5963 8897
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 6086 8888 6092 8900
rect 5951 8860 6092 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 6086 8848 6092 8860
rect 6144 8888 6150 8900
rect 6840 8888 6868 8996
rect 7024 8968 7052 8996
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 6144 8860 6868 8888
rect 6932 8888 6960 8919
rect 7006 8916 7012 8968
rect 7064 8916 7070 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 7392 8956 7420 9064
rect 7331 8928 7420 8956
rect 7469 8959 7527 8965
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 7484 8888 7512 8919
rect 6932 8860 7052 8888
rect 6144 8848 6150 8860
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 3050 8780 3056 8832
rect 3108 8780 3114 8832
rect 6825 8823 6883 8829
rect 6825 8789 6837 8823
rect 6871 8820 6883 8823
rect 6914 8820 6920 8832
rect 6871 8792 6920 8820
rect 6871 8789 6883 8792
rect 6825 8783 6883 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7024 8820 7052 8860
rect 7300 8860 7512 8888
rect 7300 8832 7328 8860
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 7024 8792 7205 8820
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 7282 8780 7288 8832
rect 7340 8780 7346 8832
rect 8128 8820 8156 8919
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8496 8900 8524 9064
rect 8757 9061 8769 9095
rect 8803 9061 8815 9095
rect 9582 9092 9588 9104
rect 8757 9055 8815 9061
rect 9048 9064 9588 9092
rect 8772 9024 8800 9055
rect 8772 8996 8984 9024
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8619 8928 8892 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8386 8848 8392 8900
rect 8444 8848 8450 8900
rect 8478 8848 8484 8900
rect 8536 8848 8542 8900
rect 8662 8820 8668 8832
rect 8128 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 8864 8820 8892 8928
rect 8956 8888 8984 8996
rect 9048 8965 9076 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 9309 9027 9367 9033
rect 9309 9024 9321 9027
rect 9140 8996 9321 9024
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9140 8888 9168 8996
rect 9309 8993 9321 8996
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9024 9459 9027
rect 9674 9024 9680 9036
rect 9447 8996 9680 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9876 9033 9904 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 11241 9095 11299 9101
rect 11241 9061 11253 9095
rect 11287 9061 11299 9095
rect 11241 9055 11299 9061
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 8956 8860 9168 8888
rect 9232 8888 9260 8919
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 9548 8928 9597 8956
rect 9548 8916 9554 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9950 8956 9956 8968
rect 9585 8919 9643 8925
rect 9692 8928 9956 8956
rect 9692 8888 9720 8928
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10594 8916 10600 8968
rect 10652 8916 10658 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11256 8956 11284 9055
rect 11422 9052 11428 9104
rect 11480 9092 11486 9104
rect 11517 9095 11575 9101
rect 11517 9092 11529 9095
rect 11480 9064 11529 9092
rect 11480 9052 11486 9064
rect 11517 9061 11529 9064
rect 11563 9061 11575 9095
rect 11517 9055 11575 9061
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 12345 9095 12403 9101
rect 12345 9092 12357 9095
rect 12216 9064 12357 9092
rect 12216 9052 12222 9064
rect 12345 9061 12357 9064
rect 12391 9061 12403 9095
rect 13354 9092 13360 9104
rect 12345 9055 12403 9061
rect 12820 9064 13360 9092
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10744 8928 11345 8956
rect 10744 8916 10750 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 9232 8860 9720 8888
rect 9769 8891 9827 8897
rect 9769 8857 9781 8891
rect 9815 8888 9827 8891
rect 10106 8891 10164 8897
rect 10106 8888 10118 8891
rect 9815 8860 10118 8888
rect 9815 8857 9827 8860
rect 9769 8851 9827 8857
rect 10106 8857 10118 8860
rect 10152 8857 10164 8891
rect 10106 8851 10164 8857
rect 9950 8820 9956 8832
rect 8864 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8820 10014 8832
rect 10612 8820 10640 8916
rect 12360 8832 12388 8919
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 12820 8965 12848 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12584 8928 12817 8956
rect 12584 8916 12590 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 12618 8848 12624 8900
rect 12676 8888 12682 8900
rect 13096 8888 13124 8919
rect 12676 8860 13124 8888
rect 12676 8848 12682 8860
rect 10008 8792 10640 8820
rect 10008 8780 10014 8792
rect 12342 8780 12348 8832
rect 12400 8780 12406 8832
rect 1104 8730 14536 8752
rect 1104 8678 4918 8730
rect 4970 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 5238 8730
rect 5290 8678 10918 8730
rect 10970 8678 10982 8730
rect 11034 8678 11046 8730
rect 11098 8678 11110 8730
rect 11162 8678 11174 8730
rect 11226 8678 11238 8730
rect 11290 8678 14536 8730
rect 1104 8656 14536 8678
rect 2498 8576 2504 8628
rect 2556 8576 2562 8628
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3326 8616 3332 8628
rect 3108 8588 3332 8616
rect 3108 8576 3114 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4798 8576 4804 8628
rect 4856 8576 4862 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6052 8588 9628 8616
rect 6052 8576 6058 8588
rect 2516 8489 2544 8576
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 4338 8548 4344 8560
rect 3016 8520 4344 8548
rect 3016 8508 3022 8520
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4816 8548 4844 8576
rect 6730 8548 6736 8560
rect 4816 8520 5856 8548
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 5828 8489 5856 8520
rect 6380 8520 6736 8548
rect 6380 8489 6408 8520
rect 6730 8508 6736 8520
rect 6788 8548 6794 8560
rect 9600 8548 9628 8588
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9824 8588 10057 8616
rect 9824 8576 9830 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 12250 8616 12256 8628
rect 12207 8588 12256 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 6788 8520 8432 8548
rect 9600 8520 9720 8548
rect 6788 8508 6794 8520
rect 8404 8492 8432 8520
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 7282 8480 7288 8492
rect 6595 8452 7288 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 5828 8412 5856 8443
rect 6178 8412 6184 8424
rect 5828 8384 6184 8412
rect 6178 8372 6184 8384
rect 6236 8412 6242 8424
rect 6564 8412 6592 8443
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 9692 8489 9720 8520
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9723 8452 9812 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 6236 8384 6592 8412
rect 6236 8372 6242 8384
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 6880 8384 7849 8412
rect 6880 8372 6886 8384
rect 7837 8381 7849 8384
rect 7883 8412 7895 8415
rect 9784 8412 9812 8452
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10060 8480 10088 8579
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 10134 8508 10140 8560
rect 10192 8548 10198 8560
rect 11698 8548 11704 8560
rect 10192 8520 11704 8548
rect 10192 8508 10198 8520
rect 11698 8508 11704 8520
rect 11756 8548 11762 8560
rect 11756 8520 12756 8548
rect 11756 8508 11762 8520
rect 12342 8480 12348 8492
rect 10060 8452 12348 8480
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 12728 8489 12756 8520
rect 13354 8508 13360 8560
rect 13412 8508 13418 8560
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13372 8480 13400 8508
rect 13127 8452 13400 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 11054 8412 11060 8424
rect 7883 8384 9720 8412
rect 9784 8384 11060 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 9692 8344 9720 8384
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 11606 8412 11612 8424
rect 11112 8384 11612 8412
rect 11112 8372 11118 8384
rect 11606 8372 11612 8384
rect 11664 8412 11670 8424
rect 11664 8384 12434 8412
rect 11664 8372 11670 8384
rect 11330 8344 11336 8356
rect 9692 8316 11336 8344
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12406 8344 12434 8384
rect 12912 8344 12940 8443
rect 12406 8316 12940 8344
rect 2314 8236 2320 8288
rect 2372 8236 2378 8288
rect 5442 8236 5448 8288
rect 5500 8236 5506 8288
rect 5813 8279 5871 8285
rect 5813 8245 5825 8279
rect 5859 8276 5871 8279
rect 6086 8276 6092 8288
rect 5859 8248 6092 8276
rect 5859 8245 5871 8248
rect 5813 8239 5871 8245
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6546 8236 6552 8288
rect 6604 8236 6610 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9677 8279 9735 8285
rect 9677 8276 9689 8279
rect 9088 8248 9689 8276
rect 9088 8236 9094 8248
rect 9677 8245 9689 8248
rect 9723 8245 9735 8279
rect 9677 8239 9735 8245
rect 1104 8186 14536 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13918 8186
rect 13970 8134 13982 8186
rect 14034 8134 14046 8186
rect 14098 8134 14110 8186
rect 14162 8134 14174 8186
rect 14226 8134 14238 8186
rect 14290 8134 14536 8186
rect 1104 8112 14536 8134
rect 4154 8032 4160 8084
rect 4212 8032 4218 8084
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4580 8044 4629 8072
rect 4580 8032 4586 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 5994 8072 6000 8084
rect 4617 8035 4675 8041
rect 4816 8044 6000 8072
rect 1486 7896 1492 7948
rect 1544 7936 1550 7948
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 1544 7908 2053 7936
rect 1544 7896 1550 7908
rect 2041 7905 2053 7908
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 3344 7908 3924 7936
rect 2056 7868 2084 7899
rect 3344 7880 3372 7908
rect 2590 7868 2596 7880
rect 2056 7840 2596 7868
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 3896 7877 3924 7908
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4706 7868 4712 7880
rect 4295 7840 4712 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4816 7877 4844 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6604 8044 6653 8072
rect 6604 8032 6610 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7374 8072 7380 8084
rect 7331 8044 7380 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8662 8032 8668 8084
rect 8720 8032 8726 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9858 8072 9864 8084
rect 9364 8044 9864 8072
rect 9364 8032 9370 8044
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10376 8044 11192 8072
rect 10376 8032 10382 8044
rect 5534 8004 5540 8016
rect 5000 7976 5540 8004
rect 5000 7877 5028 7976
rect 5534 7964 5540 7976
rect 5592 8004 5598 8016
rect 6178 8004 6184 8016
rect 5592 7976 6184 8004
rect 5592 7964 5598 7976
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 6472 7976 8953 8004
rect 5328 7939 5386 7945
rect 5328 7905 5340 7939
rect 5374 7936 5386 7939
rect 5442 7936 5448 7948
rect 5374 7908 5448 7936
rect 5374 7905 5386 7908
rect 5328 7899 5386 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 6472 7936 6500 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 9398 7964 9404 8016
rect 9456 7964 9462 8016
rect 10226 7964 10232 8016
rect 10284 7964 10290 8016
rect 11054 7964 11060 8016
rect 11112 7964 11118 8016
rect 5736 7908 6500 7936
rect 6825 7939 6883 7945
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5736 7868 5764 7908
rect 6104 7877 6132 7908
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 6914 7936 6920 7948
rect 6871 7908 6920 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 7190 7936 7196 7948
rect 6972 7908 7196 7936
rect 6972 7896 6978 7908
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7340 7908 7389 7936
rect 7340 7896 7346 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 9416 7936 9444 7964
rect 7377 7899 7435 7905
rect 7760 7908 9444 7936
rect 10244 7936 10272 7964
rect 10244 7908 10364 7936
rect 5123 7840 5764 7868
rect 5813 7871 5871 7877
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 5859 7840 5917 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5905 7837 5917 7840
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6178 7828 6184 7880
rect 6236 7828 6242 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 7006 7868 7012 7880
rect 6595 7840 7012 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 2314 7809 2320 7812
rect 2308 7800 2320 7809
rect 2275 7772 2320 7800
rect 2308 7763 2320 7772
rect 2314 7760 2320 7763
rect 2372 7760 2378 7812
rect 3800 7800 3828 7828
rect 5445 7803 5503 7809
rect 3800 7772 5212 7800
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3878 7732 3884 7744
rect 3467 7704 3884 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 4062 7732 4068 7744
rect 4019 7704 4068 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 5184 7741 5212 7772
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 5491 7772 6837 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 6932 7800 6960 7840
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 7760 7877 7788 7908
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8478 7868 8484 7880
rect 8435 7840 8484 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 7760 7800 7788 7831
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9088 7840 9413 7868
rect 9088 7828 9094 7840
rect 9401 7837 9413 7840
rect 9447 7868 9459 7871
rect 9674 7868 9680 7880
rect 9447 7840 9680 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10336 7877 10364 7908
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10597 7871 10655 7877
rect 10597 7868 10609 7871
rect 10367 7840 10609 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10597 7837 10609 7840
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 6932 7772 7788 7800
rect 8665 7803 8723 7809
rect 6825 7763 6883 7769
rect 8665 7769 8677 7803
rect 8711 7769 8723 7803
rect 8665 7763 8723 7769
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7701 5227 7735
rect 5169 7695 5227 7701
rect 5537 7735 5595 7741
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5626 7732 5632 7744
rect 5583 7704 5632 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5626 7692 5632 7704
rect 5684 7732 5690 7744
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 5684 7704 7021 7732
rect 5684 7692 5690 7704
rect 7009 7701 7021 7704
rect 7055 7701 7067 7735
rect 7009 7695 7067 7701
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7834 7732 7840 7744
rect 7699 7704 7840 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 8444 7704 8493 7732
rect 8444 7692 8450 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8680 7732 8708 7763
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 9861 7803 9919 7809
rect 9861 7800 9873 7803
rect 9640 7772 9873 7800
rect 9640 7760 9646 7772
rect 9861 7769 9873 7772
rect 9907 7769 9919 7803
rect 10244 7800 10272 7831
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 11164 7877 11192 8044
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11940 7840 11989 7868
rect 11940 7828 11946 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 10704 7800 10732 7828
rect 10244 7772 10732 7800
rect 9861 7763 9919 7769
rect 10134 7732 10140 7744
rect 8680 7704 10140 7732
rect 8481 7695 8539 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 1104 7642 14536 7664
rect 1104 7590 4918 7642
rect 4970 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 5238 7642
rect 5290 7590 10918 7642
rect 10970 7590 10982 7642
rect 11034 7590 11046 7642
rect 11098 7590 11110 7642
rect 11162 7590 11174 7642
rect 11226 7590 11238 7642
rect 11290 7590 14536 7642
rect 1104 7568 14536 7590
rect 3326 7488 3332 7540
rect 3384 7488 3390 7540
rect 3611 7531 3669 7537
rect 3611 7497 3623 7531
rect 3657 7528 3669 7531
rect 4154 7528 4160 7540
rect 3657 7500 4160 7528
rect 3657 7497 3669 7500
rect 3611 7491 3669 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5534 7528 5540 7540
rect 5399 7500 5540 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 7006 7528 7012 7540
rect 5644 7500 7012 7528
rect 3344 7460 3372 7488
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 3344 7432 3709 7460
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 3697 7423 3755 7429
rect 3786 7420 3792 7472
rect 3844 7420 3850 7472
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3476 7364 3525 7392
rect 3476 7352 3482 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3804 7391 3832 7420
rect 5261 7395 5319 7401
rect 3513 7355 3571 7361
rect 3789 7385 3847 7391
rect 3789 7351 3801 7385
rect 3835 7351 3847 7385
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5644 7392 5672 7500
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 8680 7500 10272 7528
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 7098 7460 7104 7472
rect 6144 7432 7104 7460
rect 6144 7420 6150 7432
rect 7098 7420 7104 7432
rect 7156 7460 7162 7472
rect 7469 7463 7527 7469
rect 7469 7460 7481 7463
rect 7156 7432 7481 7460
rect 7156 7420 7162 7432
rect 7469 7429 7481 7432
rect 7515 7429 7527 7463
rect 8680 7460 8708 7500
rect 10244 7472 10272 7500
rect 10502 7488 10508 7540
rect 10560 7488 10566 7540
rect 9490 7460 9496 7472
rect 7469 7423 7527 7429
rect 7852 7432 8708 7460
rect 5491 7364 5672 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 3789 7345 3847 7351
rect 5276 7324 5304 7355
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6454 7392 6460 7404
rect 6052 7364 6460 7392
rect 6052 7352 6058 7364
rect 6454 7352 6460 7364
rect 6512 7392 6518 7404
rect 6730 7392 6736 7404
rect 6512 7364 6736 7392
rect 6512 7352 6518 7364
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 5810 7324 5816 7336
rect 5276 7296 5816 7324
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 7852 7333 7880 7432
rect 8680 7401 8708 7432
rect 9140 7432 9496 7460
rect 9140 7401 9168 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 9950 7420 9956 7472
rect 10008 7420 10014 7472
rect 10226 7420 10232 7472
rect 10284 7420 10290 7472
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8665 7395 8723 7401
rect 8343 7364 8616 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7800 7296 7849 7324
rect 7800 7284 7806 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 8588 7324 8616 7364
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9125 7355 9183 7361
rect 9324 7364 9597 7392
rect 8864 7324 8892 7355
rect 9324 7336 9352 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 8588 7296 8892 7324
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 6454 7256 6460 7268
rect 3936 7228 6460 7256
rect 3936 7216 3942 7228
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 7484 7228 8769 7256
rect 7484 7200 7512 7228
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 8864 7256 8892 7296
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9548 7296 9873 7324
rect 9548 7284 9554 7296
rect 9861 7293 9873 7296
rect 9907 7324 9919 7327
rect 9968 7324 9996 7420
rect 10520 7392 10548 7488
rect 11330 7420 11336 7472
rect 11388 7460 11394 7472
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 11388 7432 11529 7460
rect 11388 7420 11394 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 11517 7423 11575 7429
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10520 7364 10609 7392
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 9907 7296 9996 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 10686 7256 10692 7268
rect 8864 7228 10692 7256
rect 8757 7219 8815 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 5718 7188 5724 7200
rect 4120 7160 5724 7188
rect 4120 7148 4126 7160
rect 5718 7148 5724 7160
rect 5776 7188 5782 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5776 7160 5825 7188
rect 5776 7148 5782 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 7892 7160 7941 7188
rect 7892 7148 7898 7160
rect 7929 7157 7941 7160
rect 7975 7188 7987 7191
rect 8570 7188 8576 7200
rect 7975 7160 8576 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 10042 7188 10048 7200
rect 9815 7160 10048 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10192 7160 10425 7188
rect 10192 7148 10198 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11790 7188 11796 7200
rect 11112 7160 11796 7188
rect 11112 7148 11118 7160
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12676 7160 12817 7188
rect 12676 7148 12682 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 1104 7098 14536 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13918 7098
rect 13970 7046 13982 7098
rect 14034 7046 14046 7098
rect 14098 7046 14110 7098
rect 14162 7046 14174 7098
rect 14226 7046 14238 7098
rect 14290 7046 14536 7098
rect 1104 7024 14536 7046
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 4706 6984 4712 6996
rect 3476 6956 4712 6984
rect 3476 6944 3482 6956
rect 4706 6944 4712 6956
rect 4764 6984 4770 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4764 6956 5181 6984
rect 4764 6944 4770 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 7834 6984 7840 6996
rect 7331 6956 7840 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9582 6984 9588 6996
rect 8444 6956 9588 6984
rect 8444 6944 8450 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10137 6987 10195 6993
rect 10137 6984 10149 6987
rect 9916 6956 10149 6984
rect 9916 6944 9922 6956
rect 10137 6953 10149 6956
rect 10183 6984 10195 6987
rect 10318 6984 10324 6996
rect 10183 6956 10324 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 11882 6984 11888 6996
rect 11440 6956 11888 6984
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 4856 6888 5580 6916
rect 4856 6876 4862 6888
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 2648 6820 3801 6848
rect 2648 6808 2654 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4396 6752 5457 6780
rect 4396 6740 4402 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 4056 6715 4114 6721
rect 4056 6681 4068 6715
rect 4102 6712 4114 6715
rect 4246 6712 4252 6724
rect 4102 6684 4252 6712
rect 4102 6681 4114 6684
rect 4056 6675 4114 6681
rect 4246 6672 4252 6684
rect 4304 6672 4310 6724
rect 5552 6721 5580 6888
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7248 6888 7665 6916
rect 7248 6876 7254 6888
rect 7653 6885 7665 6888
rect 7699 6916 7711 6919
rect 9490 6916 9496 6928
rect 7699 6888 9496 6916
rect 7699 6885 7711 6888
rect 7653 6879 7711 6885
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 9600 6916 9628 6944
rect 10229 6919 10287 6925
rect 10229 6916 10241 6919
rect 9600 6888 10241 6916
rect 10229 6885 10241 6888
rect 10275 6916 10287 6919
rect 11072 6916 11100 6944
rect 10275 6888 11100 6916
rect 10275 6885 10287 6888
rect 10229 6879 10287 6885
rect 5609 6851 5667 6857
rect 5609 6817 5621 6851
rect 5655 6848 5667 6851
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 5655 6820 6040 6848
rect 5655 6817 5667 6820
rect 5609 6811 5667 6817
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 6012 6780 6040 6820
rect 7668 6820 9597 6848
rect 6161 6783 6219 6789
rect 6161 6780 6173 6783
rect 6012 6752 6173 6780
rect 5905 6743 5963 6749
rect 6161 6749 6173 6752
rect 6207 6749 6219 6783
rect 6161 6743 6219 6749
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5626 6712 5632 6724
rect 5583 6684 5632 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 5920 6712 5948 6743
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7668 6789 7696 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6848 9827 6851
rect 10045 6851 10103 6857
rect 9815 6820 9849 6848
rect 9815 6817 9827 6820
rect 9769 6811 9827 6817
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10091 6820 10272 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7524 6752 7665 6780
rect 7524 6740 7530 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8018 6780 8024 6792
rect 7975 6752 8024 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 5828 6684 5948 6712
rect 5828 6656 5856 6684
rect 6362 6672 6368 6724
rect 6420 6712 6426 6724
rect 6420 6684 7328 6712
rect 6420 6672 6426 6684
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5442 6644 5448 6656
rect 5399 6616 5448 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5810 6604 5816 6656
rect 5868 6604 5874 6656
rect 7300 6644 7328 6684
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 7300 6616 8953 6644
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 9140 6644 9168 6743
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 9447 6783 9505 6789
rect 9447 6749 9459 6783
rect 9493 6780 9505 6783
rect 9784 6780 9812 6811
rect 10244 6792 10272 6820
rect 9493 6752 9812 6780
rect 9493 6749 9505 6752
rect 9447 6743 9505 6749
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 9784 6712 9812 6752
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 10686 6780 10692 6792
rect 10643 6752 10692 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 10686 6740 10692 6752
rect 10744 6780 10750 6792
rect 11440 6789 11468 6956
rect 11882 6944 11888 6956
rect 11940 6984 11946 6996
rect 12250 6984 12256 6996
rect 11940 6956 12256 6984
rect 11940 6944 11946 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 11425 6783 11483 6789
rect 10744 6752 11284 6780
rect 10744 6740 10750 6752
rect 9784 6684 10824 6712
rect 10796 6656 10824 6684
rect 9766 6644 9772 6656
rect 9140 6616 9772 6644
rect 8941 6607 8999 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10778 6604 10784 6656
rect 10836 6604 10842 6656
rect 11256 6653 11284 6752
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 12618 6780 12624 6792
rect 11563 6752 12624 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 11762 6715 11820 6721
rect 11762 6712 11774 6715
rect 11388 6684 11774 6712
rect 11388 6672 11394 6684
rect 11762 6681 11774 6684
rect 11808 6681 11820 6715
rect 11762 6675 11820 6681
rect 11241 6647 11299 6653
rect 11241 6613 11253 6647
rect 11287 6644 11299 6647
rect 12158 6644 12164 6656
rect 11287 6616 12164 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12308 6616 12909 6644
rect 12308 6604 12314 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 1104 6554 14536 6576
rect 1104 6502 4918 6554
rect 4970 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 5238 6554
rect 5290 6502 10918 6554
rect 10970 6502 10982 6554
rect 11034 6502 11046 6554
rect 11098 6502 11110 6554
rect 11162 6502 11174 6554
rect 11226 6502 11238 6554
rect 11290 6502 14536 6554
rect 1104 6480 14536 6502
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 8536 6412 10180 6440
rect 8536 6400 8542 6412
rect 2216 6375 2274 6381
rect 2216 6341 2228 6375
rect 2262 6372 2274 6375
rect 2406 6372 2412 6384
rect 2262 6344 2412 6372
rect 2262 6341 2274 6344
rect 2216 6335 2274 6341
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 7742 6332 7748 6384
rect 7800 6332 7806 6384
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 8665 6375 8723 6381
rect 8665 6372 8677 6375
rect 8076 6344 8677 6372
rect 8076 6332 8082 6344
rect 8665 6341 8677 6344
rect 8711 6341 8723 6375
rect 8665 6335 8723 6341
rect 9858 6332 9864 6384
rect 9916 6332 9922 6384
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6304 4951 6307
rect 4939 6276 5396 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1728 6208 1961 6236
rect 1728 6196 1734 6208
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6236 3847 6239
rect 4062 6236 4068 6248
rect 3835 6208 4068 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 4062 6196 4068 6208
rect 4120 6236 4126 6248
rect 5166 6236 5172 6248
rect 4120 6208 5172 6236
rect 4120 6196 4126 6208
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5368 6245 5396 6276
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5767 6276 5825 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 7760 6304 7788 6332
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7760 6276 7849 6304
rect 5813 6267 5871 6273
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8386 6304 8392 6316
rect 8343 6276 8392 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5442 6236 5448 6248
rect 5399 6208 5448 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 4246 6168 4252 6180
rect 3344 6140 4252 6168
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 3344 6109 3372 6140
rect 4246 6128 4252 6140
rect 4304 6128 4310 6180
rect 8128 6168 8156 6267
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 8628 6276 8769 6304
rect 8628 6264 8634 6276
rect 8757 6273 8769 6276
rect 8803 6304 8815 6307
rect 9769 6307 9827 6313
rect 8803 6302 9674 6304
rect 9769 6302 9781 6307
rect 8803 6276 9781 6302
rect 8803 6273 8815 6276
rect 9646 6274 9781 6276
rect 8757 6267 8815 6273
rect 9769 6273 9781 6274
rect 9815 6304 9827 6307
rect 9876 6304 9904 6332
rect 10033 6317 10091 6323
rect 9815 6276 9904 6304
rect 9947 6307 10005 6313
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9947 6273 9959 6307
rect 9993 6273 10005 6307
rect 10033 6283 10045 6317
rect 10079 6283 10091 6317
rect 10033 6277 10091 6283
rect 10152 6304 10180 6412
rect 10226 6400 10232 6452
rect 10284 6400 10290 6452
rect 11050 6443 11108 6449
rect 11050 6409 11062 6443
rect 11096 6440 11108 6443
rect 11330 6440 11336 6452
rect 11096 6412 11336 6440
rect 11096 6409 11108 6412
rect 11050 6403 11108 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 13814 6440 13820 6452
rect 12544 6412 13820 6440
rect 10244 6372 10272 6400
rect 10244 6344 10640 6372
rect 10612 6313 10640 6344
rect 11701 6317 11759 6323
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9947 6267 10005 6273
rect 8128 6140 9628 6168
rect 9600 6112 9628 6140
rect 9766 6128 9772 6180
rect 9824 6128 9830 6180
rect 9968 6168 9996 6267
rect 10060 6248 10088 6277
rect 10152 6276 10241 6304
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 10686 6264 10692 6316
rect 10744 6264 10750 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10796 6276 10885 6304
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10318 6196 10324 6248
rect 10376 6196 10382 6248
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10704 6236 10732 6264
rect 10459 6208 10732 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10226 6168 10232 6180
rect 9968 6140 10232 6168
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 1636 6072 3341 6100
rect 1636 6060 1642 6072
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3329 6063 3387 6069
rect 3418 6060 3424 6112
rect 3476 6060 3482 6112
rect 5997 6103 6055 6109
rect 5997 6069 6009 6103
rect 6043 6100 6055 6103
rect 6086 6100 6092 6112
rect 6043 6072 6092 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 7653 6103 7711 6109
rect 7653 6069 7665 6103
rect 7699 6100 7711 6103
rect 7834 6100 7840 6112
rect 7699 6072 7840 6100
rect 7699 6069 7711 6072
rect 7653 6063 7711 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 10428 6100 10456 6199
rect 10796 6109 10824 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11701 6283 11713 6317
rect 11747 6283 11759 6317
rect 11701 6277 11759 6283
rect 11885 6307 11943 6313
rect 11716 6248 11744 6277
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 12253 6307 12311 6313
rect 11931 6276 12204 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 11698 6196 11704 6248
rect 11756 6196 11762 6248
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 11992 6168 12020 6199
rect 12066 6196 12072 6248
rect 12124 6196 12130 6248
rect 12176 6236 12204 6276
rect 12253 6273 12265 6307
rect 12299 6304 12311 6307
rect 12544 6304 12572 6412
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 12676 6344 13952 6372
rect 12676 6332 12682 6344
rect 13924 6313 13952 6344
rect 12299 6276 12572 6304
rect 13653 6307 13711 6313
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 13653 6273 13665 6307
rect 13699 6304 13711 6307
rect 13909 6307 13967 6313
rect 13699 6276 13860 6304
rect 13699 6273 13711 6276
rect 13653 6267 13711 6273
rect 12342 6236 12348 6248
rect 12176 6208 12348 6236
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12802 6236 12808 6248
rect 12483 6208 12808 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 13832 6236 13860 6276
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14458 6236 14464 6248
rect 13832 6208 14464 6236
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 12894 6168 12900 6180
rect 10928 6140 11744 6168
rect 11992 6140 12900 6168
rect 10928 6128 10934 6140
rect 9640 6072 10456 6100
rect 10781 6103 10839 6109
rect 9640 6060 9646 6072
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 11606 6100 11612 6112
rect 10827 6072 11612 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11716 6100 11744 6140
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 11716 6072 12541 6100
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 1104 6010 14536 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13918 6010
rect 13970 5958 13982 6010
rect 14034 5958 14046 6010
rect 14098 5958 14110 6010
rect 14162 5958 14174 6010
rect 14226 5958 14238 6010
rect 14290 5958 14536 6010
rect 1104 5936 14536 5958
rect 2406 5856 2412 5908
rect 2464 5856 2470 5908
rect 3418 5896 3424 5908
rect 2746 5868 3424 5896
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2746 5692 2774 5868
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3660 5868 3801 5896
rect 3660 5856 3666 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 5534 5896 5540 5908
rect 5031 5868 5540 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 5960 5868 8217 5896
rect 5960 5856 5966 5868
rect 8205 5865 8217 5868
rect 8251 5896 8263 5899
rect 8386 5896 8392 5908
rect 8251 5868 8392 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 9214 5896 9220 5908
rect 8711 5868 9220 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 6270 5828 6276 5840
rect 4080 5800 6276 5828
rect 4080 5701 4108 5800
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 8478 5828 8484 5840
rect 7576 5800 8484 5828
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 5224 5732 7144 5760
rect 5224 5720 5230 5732
rect 2639 5664 2774 5692
rect 3973 5695 4031 5701
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 3602 5584 3608 5636
rect 3660 5624 3666 5636
rect 3988 5624 4016 5655
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4304 5664 4353 5692
rect 4304 5652 4310 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 4341 5655 4399 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4522 5692 4528 5704
rect 4479 5664 4528 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 4847 5664 6592 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 3660 5596 4099 5624
rect 3660 5584 3666 5596
rect 4071 5556 4099 5596
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4617 5627 4675 5633
rect 4617 5624 4629 5627
rect 4212 5596 4629 5624
rect 4212 5584 4218 5596
rect 4617 5593 4629 5596
rect 4663 5593 4675 5627
rect 4617 5587 4675 5593
rect 4816 5556 4844 5655
rect 6564 5636 6592 5664
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 5626 5584 5632 5636
rect 5684 5624 5690 5636
rect 5684 5596 6500 5624
rect 5684 5584 5690 5596
rect 4071 5528 4844 5556
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 5810 5556 5816 5568
rect 5583 5528 5816 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 6472 5556 6500 5596
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 6917 5627 6975 5633
rect 6917 5624 6929 5627
rect 6604 5596 6929 5624
rect 6604 5584 6610 5596
rect 6917 5593 6929 5596
rect 6963 5593 6975 5627
rect 7116 5624 7144 5732
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5692 7251 5695
rect 7576 5692 7604 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8680 5760 8708 5859
rect 9214 5856 9220 5868
rect 9272 5896 9278 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 9272 5868 9321 5896
rect 9272 5856 9278 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 10870 5896 10876 5908
rect 9456 5868 10876 5896
rect 9456 5856 9462 5868
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 11606 5856 11612 5908
rect 11664 5856 11670 5908
rect 11790 5856 11796 5908
rect 11848 5856 11854 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 12124 5868 12357 5896
rect 12124 5856 12130 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 9582 5828 9588 5840
rect 8036 5732 8708 5760
rect 9232 5800 9588 5828
rect 8036 5701 8064 5732
rect 7239 5664 7604 5692
rect 7653 5695 7711 5701
rect 7239 5661 7251 5664
rect 7193 5655 7251 5661
rect 7653 5661 7665 5695
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 7668 5624 7696 5655
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 9232 5692 9260 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 10226 5828 10232 5840
rect 9692 5800 10232 5828
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 9692 5760 9720 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 10594 5788 10600 5840
rect 10652 5788 10658 5840
rect 11164 5828 11192 5856
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 11164 5800 11713 5828
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11808 5828 11836 5856
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 11808 5800 12173 5828
rect 11701 5791 11759 5797
rect 12161 5797 12173 5800
rect 12207 5797 12219 5831
rect 12161 5791 12219 5797
rect 10042 5760 10048 5772
rect 9447 5732 9720 5760
rect 9968 5732 10048 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 8527 5664 9260 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9766 5692 9772 5704
rect 9600 5664 9772 5692
rect 7834 5624 7840 5636
rect 7116 5596 7604 5624
rect 7668 5596 7840 5624
rect 6917 5587 6975 5593
rect 7098 5556 7104 5568
rect 6472 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7576 5556 7604 5596
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 9600 5556 9628 5664
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 9968 5701 9996 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10612 5760 10640 5788
rect 11793 5763 11851 5769
rect 10192 5732 10640 5760
rect 11256 5732 11652 5760
rect 10192 5720 10198 5732
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 9692 5596 9873 5624
rect 9692 5565 9720 5596
rect 9861 5593 9873 5596
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 7576 5528 9628 5556
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5525 9735 5559
rect 10244 5556 10272 5655
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 11256 5701 11284 5732
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 10836 5664 11253 5692
rect 10836 5652 10842 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11422 5652 11428 5704
rect 11480 5652 11486 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 11624 5692 11652 5732
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 12066 5760 12072 5772
rect 11839 5732 12072 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 11808 5692 11928 5694
rect 12342 5692 12348 5704
rect 11624 5666 12348 5692
rect 11624 5664 11836 5666
rect 11900 5664 12348 5666
rect 11517 5655 11575 5661
rect 10321 5627 10379 5633
rect 10321 5593 10333 5627
rect 10367 5624 10379 5627
rect 10502 5624 10508 5636
rect 10367 5596 10508 5624
rect 10367 5593 10379 5596
rect 10321 5587 10379 5593
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 10962 5624 10968 5636
rect 10652 5596 10968 5624
rect 10652 5584 10658 5596
rect 10962 5584 10968 5596
rect 11020 5624 11026 5636
rect 11532 5624 11560 5655
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12618 5692 12624 5704
rect 12575 5664 12624 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 12802 5701 12808 5704
rect 12796 5692 12808 5701
rect 12763 5664 12808 5692
rect 12796 5655 12808 5664
rect 12802 5652 12808 5655
rect 12860 5652 12866 5704
rect 11020 5596 11560 5624
rect 11020 5584 11026 5596
rect 11882 5584 11888 5636
rect 11940 5584 11946 5636
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 13538 5624 13544 5636
rect 12032 5596 13544 5624
rect 12032 5584 12038 5596
rect 13538 5584 13544 5596
rect 13596 5584 13602 5636
rect 10778 5556 10784 5568
rect 10244 5528 10784 5556
rect 9677 5519 9735 5525
rect 10778 5516 10784 5528
rect 10836 5556 10842 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10836 5528 11345 5556
rect 10836 5516 10842 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 11992 5556 12020 5584
rect 11480 5528 12020 5556
rect 11480 5516 11486 5528
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 13909 5559 13967 5565
rect 13909 5556 13921 5559
rect 13872 5528 13921 5556
rect 13872 5516 13878 5528
rect 13909 5525 13921 5528
rect 13955 5556 13967 5559
rect 14550 5556 14556 5568
rect 13955 5528 14556 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 1104 5466 14536 5488
rect 1104 5414 4918 5466
rect 4970 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 5238 5466
rect 5290 5414 10918 5466
rect 10970 5414 10982 5466
rect 11034 5414 11046 5466
rect 11098 5414 11110 5466
rect 11162 5414 11174 5466
rect 11226 5414 11238 5466
rect 11290 5414 14536 5466
rect 1104 5392 14536 5414
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 3513 5287 3571 5293
rect 3513 5253 3525 5287
rect 3559 5253 3571 5287
rect 3513 5247 3571 5253
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 2372 5188 3249 5216
rect 2372 5176 2378 5188
rect 3237 5185 3249 5188
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3436 5080 3464 5179
rect 3528 5148 3556 5247
rect 3602 5176 3608 5228
rect 3660 5176 3666 5228
rect 3804 5216 3832 5315
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4580 5324 4813 5352
rect 4580 5312 4586 5324
rect 4801 5321 4813 5324
rect 4847 5352 4859 5355
rect 8754 5352 8760 5364
rect 4847 5324 8760 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 9306 5352 9312 5364
rect 9079 5324 9312 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9490 5312 9496 5364
rect 9548 5312 9554 5364
rect 11790 5312 11796 5364
rect 11848 5312 11854 5364
rect 12710 5352 12716 5364
rect 12406 5324 12716 5352
rect 6086 5244 6092 5296
rect 6144 5244 6150 5296
rect 8294 5284 8300 5296
rect 7668 5256 8300 5284
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3804 5188 4077 5216
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4430 5216 4436 5228
rect 4065 5179 4123 5185
rect 4172 5188 4436 5216
rect 4172 5148 4200 5188
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 5925 5219 5983 5225
rect 5925 5185 5937 5219
rect 5971 5216 5983 5219
rect 6104 5216 6132 5244
rect 5971 5188 6132 5216
rect 5971 5185 5983 5188
rect 5925 5179 5983 5185
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7668 5225 7696 5256
rect 8294 5244 8300 5256
rect 8352 5284 8358 5296
rect 9508 5284 9536 5312
rect 8352 5256 9536 5284
rect 8352 5244 8358 5256
rect 8956 5225 8984 5256
rect 10410 5244 10416 5296
rect 10468 5284 10474 5296
rect 10468 5256 10916 5284
rect 10468 5244 10474 5256
rect 7653 5219 7711 5225
rect 6788 5188 7604 5216
rect 6788 5176 6794 5188
rect 3528 5120 4200 5148
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5117 6239 5151
rect 6564 5148 6592 5176
rect 6822 5148 6828 5160
rect 6564 5120 6828 5148
rect 6181 5111 6239 5117
rect 4154 5080 4160 5092
rect 3436 5052 4160 5080
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3384 4984 3893 5012
rect 3384 4972 3390 4984
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4264 5012 4292 5111
rect 4120 4984 4292 5012
rect 4120 4972 4126 4984
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6196 5012 6224 5111
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 6457 5083 6515 5089
rect 6457 5049 6469 5083
rect 6503 5080 6515 5083
rect 7576 5080 7604 5188
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9582 5216 9588 5228
rect 9171 5188 9588 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 9140 5148 9168 5179
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 10778 5216 10784 5228
rect 10735 5188 10784 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 10888 5225 10916 5256
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 10962 5216 10968 5228
rect 10919 5188 10968 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11808 5216 11836 5312
rect 12406 5284 12434 5324
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 13630 5312 13636 5364
rect 13688 5312 13694 5364
rect 11992 5256 12434 5284
rect 12912 5284 12940 5312
rect 12912 5256 13216 5284
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11808 5188 11897 5216
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 7975 5120 9168 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 11992 5080 12020 5256
rect 13188 5228 13216 5256
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12400 5188 12909 5216
rect 12400 5176 12406 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13170 5176 13176 5228
rect 13228 5176 13234 5228
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13556 5148 13584 5179
rect 13814 5176 13820 5228
rect 13872 5176 13878 5228
rect 12768 5120 13584 5148
rect 12768 5108 12774 5120
rect 6503 5052 6684 5080
rect 7576 5052 12020 5080
rect 6503 5049 6515 5052
rect 6457 5043 6515 5049
rect 6656 5024 6684 5052
rect 5868 4984 6224 5012
rect 5868 4972 5874 4984
rect 6638 4972 6644 5024
rect 6696 4972 6702 5024
rect 7834 4972 7840 5024
rect 7892 4972 7898 5024
rect 8205 5015 8263 5021
rect 8205 4981 8217 5015
rect 8251 5012 8263 5015
rect 8386 5012 8392 5024
rect 8251 4984 8392 5012
rect 8251 4981 8263 4984
rect 8205 4975 8263 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 10686 4972 10692 5024
rect 10744 4972 10750 5024
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11020 4984 11989 5012
rect 11020 4972 11026 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 11977 4975 12035 4981
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 12308 4984 12449 5012
rect 12308 4972 12314 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12437 4975 12495 4981
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14047 4984 14596 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 1104 4922 14536 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13918 4922
rect 13970 4870 13982 4922
rect 14034 4870 14046 4922
rect 14098 4870 14110 4922
rect 14162 4870 14174 4922
rect 14226 4870 14238 4922
rect 14290 4870 14536 4922
rect 1104 4848 14536 4870
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 10778 4808 10784 4820
rect 8904 4780 10784 4808
rect 8904 4768 8910 4780
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 11882 4808 11888 4820
rect 11839 4780 11888 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 14568 4808 14596 4984
rect 12299 4780 14596 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 9125 4743 9183 4749
rect 9125 4709 9137 4743
rect 9171 4740 9183 4743
rect 9306 4740 9312 4752
rect 9171 4712 9312 4740
rect 9171 4709 9183 4712
rect 9125 4703 9183 4709
rect 9306 4700 9312 4712
rect 9364 4700 9370 4752
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 3752 4644 4108 4672
rect 3752 4632 3758 4644
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 1670 4604 1676 4616
rect 1627 4576 1676 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 4080 4613 4108 4644
rect 6472 4644 8616 4672
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 1848 4539 1906 4545
rect 1848 4505 1860 4539
rect 1894 4536 1906 4539
rect 2038 4536 2044 4548
rect 1894 4508 2044 4536
rect 1894 4505 1906 4508
rect 1848 4499 1906 4505
rect 2038 4496 2044 4508
rect 2096 4496 2102 4548
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2372 4440 2973 4468
rect 2372 4428 2378 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 3988 4468 4016 4567
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 6472 4613 6500 4644
rect 8588 4616 8616 4644
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 8570 4564 8576 4616
rect 8628 4564 8634 4616
rect 9214 4604 9220 4616
rect 8680 4576 9220 4604
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 4798 4536 4804 4548
rect 4212 4508 4804 4536
rect 4212 4496 4218 4508
rect 4798 4496 4804 4508
rect 4856 4536 4862 4548
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 4856 4508 6653 4536
rect 4856 4496 4862 4508
rect 6641 4505 6653 4508
rect 6687 4536 6699 4539
rect 8496 4536 8524 4564
rect 8680 4536 8708 4576
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10336 4576 10425 4604
rect 6687 4508 6776 4536
rect 8496 4508 8708 4536
rect 6687 4505 6699 4508
rect 6641 4499 6699 4505
rect 6748 4480 6776 4508
rect 8938 4496 8944 4548
rect 8996 4496 9002 4548
rect 10336 4480 10364 4576
rect 10413 4573 10425 4576
rect 10459 4604 10471 4607
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 10459 4576 12541 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 12529 4573 12541 4576
rect 12575 4604 12587 4607
rect 12618 4604 12624 4616
rect 12575 4576 12624 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 10658 4539 10716 4545
rect 10658 4536 10670 4539
rect 10560 4508 10670 4536
rect 10560 4496 10566 4508
rect 10658 4505 10670 4508
rect 10704 4505 10716 4539
rect 10658 4499 10716 4505
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 10836 4508 12081 4536
rect 10836 4496 10842 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 12069 4499 12127 4505
rect 12250 4496 12256 4548
rect 12308 4545 12314 4548
rect 12802 4545 12808 4548
rect 12308 4539 12343 4545
rect 12331 4505 12343 4539
rect 12308 4499 12343 4505
rect 12796 4499 12808 4545
rect 12308 4496 12314 4499
rect 12802 4496 12808 4499
rect 12860 4496 12866 4548
rect 4614 4468 4620 4480
rect 3988 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 6730 4428 6736 4480
rect 6788 4428 6794 4480
rect 7006 4428 7012 4480
rect 7064 4428 7070 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8352 4440 9229 4468
rect 8352 4428 8358 4440
rect 9217 4437 9229 4440
rect 9263 4468 9275 4471
rect 9398 4468 9404 4480
rect 9263 4440 9404 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10318 4428 10324 4480
rect 10376 4428 10382 4480
rect 12434 4428 12440 4480
rect 12492 4428 12498 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 13909 4471 13967 4477
rect 13909 4468 13921 4471
rect 13872 4440 13921 4468
rect 13872 4428 13878 4440
rect 13909 4437 13921 4440
rect 13955 4468 13967 4471
rect 14366 4468 14372 4480
rect 13955 4440 14372 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 1104 4378 14536 4400
rect 1104 4326 4918 4378
rect 4970 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 5238 4378
rect 5290 4326 10918 4378
rect 10970 4326 10982 4378
rect 11034 4326 11046 4378
rect 11098 4326 11110 4378
rect 11162 4326 11174 4378
rect 11226 4326 11238 4378
rect 11290 4326 14536 4378
rect 1104 4304 14536 4326
rect 2038 4224 2044 4276
rect 2096 4224 2102 4276
rect 3786 4224 3792 4276
rect 3844 4224 3850 4276
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 5445 4267 5503 4273
rect 4028 4236 5212 4264
rect 4028 4224 4034 4236
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 3326 4128 3332 4140
rect 2271 4100 3332 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3804 4128 3832 4224
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 4798 4196 4804 4208
rect 4479 4168 4804 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 4798 4156 4804 4168
rect 4856 4196 4862 4208
rect 5184 4205 5212 4236
rect 5445 4233 5457 4267
rect 5491 4233 5503 4267
rect 6822 4264 6828 4276
rect 5445 4227 5503 4233
rect 6564 4236 6828 4264
rect 5077 4199 5135 4205
rect 5077 4196 5089 4199
rect 4856 4168 5089 4196
rect 4856 4156 4862 4168
rect 5077 4165 5089 4168
rect 5123 4165 5135 4199
rect 5077 4159 5135 4165
rect 5169 4199 5227 4205
rect 5169 4165 5181 4199
rect 5215 4165 5227 4199
rect 5169 4159 5227 4165
rect 3467 4100 3832 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 4062 4060 4068 4072
rect 3651 4032 4068 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 4540 3992 4568 4091
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 4890 4088 4896 4140
rect 4948 4088 4954 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 5000 4100 5273 4128
rect 4632 4060 4660 4088
rect 5000 4060 5028 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5460 4128 5488 4227
rect 6564 4137 6592 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7006 4224 7012 4276
rect 7064 4224 7070 4276
rect 8297 4267 8355 4273
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8938 4264 8944 4276
rect 8343 4236 8944 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9306 4224 9312 4276
rect 9364 4224 9370 4276
rect 9766 4224 9772 4276
rect 9824 4224 9830 4276
rect 12434 4224 12440 4276
rect 12492 4224 12498 4276
rect 12802 4224 12808 4276
rect 12860 4224 12866 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13228 4236 13645 4264
rect 13228 4224 13234 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 6730 4156 6736 4208
rect 6788 4156 6794 4208
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5460 4100 5733 4128
rect 5261 4091 5319 4097
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 5721 4091 5779 4097
rect 5828 4100 6561 4128
rect 4632 4032 5028 4060
rect 5276 4060 5304 4091
rect 5828 4060 5856 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6638 4088 6644 4140
rect 6696 4088 6702 4140
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 7024 4128 7052 4224
rect 8386 4156 8392 4208
rect 8444 4156 8450 4208
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7024 4100 7205 4128
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8294 4128 8300 4140
rect 8159 4100 8300 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9030 4088 9036 4140
rect 9088 4088 9094 4140
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 9324 4137 9352 4224
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 9674 4196 9680 4208
rect 9456 4168 9680 4196
rect 9456 4156 9462 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 9784 4159 9812 4224
rect 9766 4153 9824 4159
rect 9858 4156 9864 4208
rect 9916 4156 9922 4208
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9766 4119 9778 4153
rect 9812 4119 9824 4153
rect 9766 4113 9824 4119
rect 10045 4131 10103 4137
rect 9585 4091 9643 4097
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10091 4100 10548 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 5276 4032 5856 4060
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 3200 3964 4568 3992
rect 3200 3952 3206 3964
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 5920 3992 5948 4023
rect 7024 3992 7052 4023
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7156 4032 8033 4060
rect 7156 4020 7162 4032
rect 8021 4029 8033 4032
rect 8067 4060 8079 4063
rect 9122 4060 9128 4072
rect 8067 4032 9128 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9232 4060 9260 4088
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 9232 4032 9413 4060
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9600 4060 9628 4091
rect 10520 4072 10548 4100
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10744 4100 10793 4128
rect 10744 4088 10750 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 12452 4128 12480 4224
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12452 4100 12633 4128
rect 10781 4091 10839 4097
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 9858 4060 9864 4072
rect 9600 4032 9864 4060
rect 9401 4023 9459 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 10502 4020 10508 4072
rect 10560 4020 10566 4072
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10652 4032 10977 4060
rect 10652 4020 10658 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 8846 3992 8852 4004
rect 5500 3964 8852 3992
rect 5500 3952 5506 3964
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3992 9551 3995
rect 9766 3992 9772 4004
rect 9539 3964 9772 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 3234 3884 3240 3936
rect 3292 3884 3298 3936
rect 4798 3884 4804 3936
rect 4856 3884 4862 3936
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 6362 3884 6368 3936
rect 6420 3884 6426 3936
rect 7374 3884 7380 3936
rect 7432 3884 7438 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7892 3896 7941 3924
rect 7892 3884 7898 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10100 3896 10241 3924
rect 10100 3884 10106 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 1104 3834 14536 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13918 3834
rect 13970 3782 13982 3834
rect 14034 3782 14046 3834
rect 14098 3782 14110 3834
rect 14162 3782 14174 3834
rect 14226 3782 14238 3834
rect 14290 3782 14536 3834
rect 1104 3760 14536 3782
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 4798 3680 4804 3732
rect 4856 3680 4862 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 5626 3720 5632 3732
rect 4948 3692 5632 3720
rect 4948 3680 4954 3692
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 6362 3720 6368 3732
rect 5736 3692 6368 3720
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 3252 3516 3280 3680
rect 4816 3584 4844 3680
rect 4632 3556 4844 3584
rect 4632 3525 4660 3556
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 5537 3587 5595 3593
rect 5537 3584 5549 3587
rect 5500 3556 5549 3584
rect 5500 3544 5506 3556
rect 5537 3553 5549 3556
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 2915 3488 3280 3516
rect 4617 3519 4675 3525
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 5460 3516 5488 3544
rect 5736 3525 5764 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7374 3680 7380 3732
rect 7432 3680 7438 3732
rect 9766 3680 9772 3732
rect 9824 3680 9830 3732
rect 4847 3488 5488 3516
rect 5721 3519 5779 3525
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 5721 3485 5733 3519
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5868 3488 6009 3516
rect 5868 3476 5874 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 7392 3516 7420 3680
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 7392 3488 7665 3516
rect 5997 3479 6055 3485
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9088 3488 9505 3516
rect 9088 3476 9094 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 10502 3516 10508 3528
rect 9631 3488 10508 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 6264 3451 6322 3457
rect 6264 3417 6276 3451
rect 6310 3448 6322 3451
rect 6362 3448 6368 3460
rect 6310 3420 6368 3448
rect 6310 3417 6322 3420
rect 6264 3411 6322 3417
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 8404 3448 8432 3476
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 8404 3420 9781 3448
rect 9769 3417 9781 3420
rect 9815 3448 9827 3451
rect 10594 3448 10600 3460
rect 9815 3420 10600 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 2682 3340 2688 3392
rect 2740 3340 2746 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 4212 3352 4445 3380
rect 4212 3340 4218 3352
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 4433 3343 4491 3349
rect 5902 3340 5908 3392
rect 5960 3340 5966 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7377 3383 7435 3389
rect 7377 3380 7389 3383
rect 6972 3352 7389 3380
rect 6972 3340 6978 3352
rect 7377 3349 7389 3352
rect 7423 3349 7435 3383
rect 7377 3343 7435 3349
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 1104 3290 14536 3312
rect 1104 3238 4918 3290
rect 4970 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 5238 3290
rect 5290 3238 10918 3290
rect 10970 3238 10982 3290
rect 11034 3238 11046 3290
rect 11098 3238 11110 3290
rect 11162 3238 11174 3290
rect 11226 3238 11238 3290
rect 11290 3238 14536 3290
rect 1104 3216 14536 3238
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4304 3148 4537 3176
rect 4304 3136 4310 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 5994 3176 6000 3188
rect 5684 3148 6000 3176
rect 5684 3136 5690 3148
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6362 3136 6368 3188
rect 6420 3136 6426 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 9088 3148 9137 3176
rect 9088 3136 9094 3148
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9125 3139 9183 3145
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 14001 3179 14059 3185
rect 14001 3145 14013 3179
rect 14047 3176 14059 3179
rect 14458 3176 14464 3188
rect 14047 3148 14464 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 5810 3108 5816 3120
rect 3160 3080 5816 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 3160 3049 3188 3080
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 1728 3012 3157 3040
rect 1728 3000 1734 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3412 3043 3470 3049
rect 3412 3009 3424 3043
rect 3458 3040 3470 3043
rect 3786 3040 3792 3052
rect 3458 3012 3792 3040
rect 3458 3009 3470 3012
rect 3412 3003 3470 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4632 3049 4660 3080
rect 5810 3068 5816 3080
rect 5868 3108 5874 3120
rect 7098 3108 7104 3120
rect 5868 3080 7104 3108
rect 5868 3068 5874 3080
rect 7098 3068 7104 3080
rect 7156 3108 7162 3120
rect 7156 3080 7788 3108
rect 7156 3068 7162 3080
rect 4890 3049 4896 3052
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4884 3003 4896 3049
rect 4890 3000 4896 3003
rect 4948 3000 4954 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 7760 3049 7788 3080
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 7990 3111 8048 3117
rect 7990 3108 8002 3111
rect 7892 3080 8002 3108
rect 7892 3068 7898 3080
rect 7990 3077 8002 3080
rect 8036 3077 8048 3111
rect 7990 3071 8048 3077
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5960 3012 6561 3040
rect 5960 3000 5966 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 10428 3040 10456 3136
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10428 3012 10701 3040
rect 7745 3003 7803 3009
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 12888 3043 12946 3049
rect 12888 3009 12900 3043
rect 12934 3040 12946 3043
rect 13446 3040 13452 3052
rect 12934 3012 13452 3040
rect 12934 3009 12946 3012
rect 12888 3003 12946 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2836 10931 2839
rect 11054 2836 11060 2848
rect 10919 2808 11060 2836
rect 10919 2805 10931 2808
rect 10873 2799 10931 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 1104 2746 14536 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13918 2746
rect 13970 2694 13982 2746
rect 14034 2694 14046 2746
rect 14098 2694 14110 2746
rect 14162 2694 14174 2746
rect 14226 2694 14238 2746
rect 14290 2694 14536 2746
rect 1104 2672 14536 2694
rect 3786 2592 3792 2644
rect 3844 2592 3850 2644
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4304 2604 4568 2632
rect 4304 2592 4310 2604
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2564 3663 2567
rect 3651 2536 4292 2564
rect 3651 2533 3663 2536
rect 3605 2527 3663 2533
rect 1670 2456 1676 2508
rect 1728 2496 1734 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1728 2468 2237 2496
rect 1728 2456 1734 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2314 2428 2320 2440
rect 2179 2400 2320 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2498 2437 2504 2440
rect 2492 2428 2504 2437
rect 2459 2400 2504 2428
rect 2492 2391 2504 2400
rect 2498 2388 2504 2391
rect 2556 2388 2562 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4154 2428 4160 2440
rect 4019 2400 4160 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 4264 2437 4292 2536
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4338 2428 4344 2440
rect 4295 2400 4344 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4540 2428 4568 2604
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4948 2604 4997 2632
rect 4948 2592 4954 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8628 2604 10456 2632
rect 8628 2592 8634 2604
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 7156 2468 7205 2496
rect 7156 2456 7162 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4540 2400 4905 2428
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5626 2428 5632 2440
rect 5215 2400 5632 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 6052 2400 6193 2428
rect 6052 2388 6058 2400
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7466 2437 7472 2440
rect 7460 2428 7472 2437
rect 7427 2400 7472 2428
rect 7460 2391 7472 2400
rect 7466 2388 7472 2391
rect 7524 2388 7530 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10318 2428 10324 2440
rect 9263 2400 10324 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10428 2428 10456 2604
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10560 2604 10609 2632
rect 10560 2592 10566 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 13446 2592 13452 2644
rect 13504 2592 13510 2644
rect 11054 2456 11060 2508
rect 11112 2456 11118 2508
rect 14366 2496 14372 2508
rect 12636 2468 14372 2496
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10428 2400 10885 2428
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 11072 2428 11100 2456
rect 12636 2437 12664 2468
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11072 2400 11345 2428
rect 10873 2391 10931 2397
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2428 13967 2431
rect 14458 2428 14464 2440
rect 13955 2400 14464 2428
rect 13955 2397 13967 2400
rect 13909 2391 13967 2397
rect 9306 2320 9312 2372
rect 9364 2360 9370 2372
rect 9462 2363 9520 2369
rect 9462 2360 9474 2363
rect 9364 2332 9474 2360
rect 9364 2320 9370 2332
rect 9462 2329 9474 2332
rect 9508 2329 9520 2363
rect 9462 2323 9520 2329
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 13648 2360 13676 2391
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 14918 2360 14924 2372
rect 9824 2332 10732 2360
rect 13648 2332 14924 2360
rect 9824 2320 9830 2332
rect 750 2252 756 2304
rect 808 2292 814 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 808 2264 1409 2292
rect 808 2252 814 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 1946 2252 1952 2304
rect 2004 2252 2010 2304
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3752 2264 4077 2292
rect 3752 2252 3758 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 5994 2252 6000 2304
rect 6052 2252 6058 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 10704 2301 10732 2332
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 8720 2264 8953 2292
rect 8720 2252 8726 2264
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 8941 2255 8999 2261
rect 10689 2295 10747 2301
rect 10689 2261 10701 2295
rect 10735 2261 10747 2295
rect 10689 2255 10747 2261
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11330 2292 11336 2304
rect 11195 2264 11336 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11330 2252 11336 2264
rect 11388 2252 11394 2304
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12400 2264 12449 2292
rect 12400 2252 12406 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 13722 2252 13728 2304
rect 13780 2252 13786 2304
rect 1104 2202 14536 2224
rect 1104 2150 4918 2202
rect 4970 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 5238 2202
rect 5290 2150 10918 2202
rect 10970 2150 10982 2202
rect 11034 2150 11046 2202
rect 11098 2150 11110 2202
rect 11162 2150 11174 2202
rect 11226 2150 11238 2202
rect 11290 2150 14536 2202
rect 1104 2128 14536 2150
<< via1 >>
rect 4918 15206 4970 15258
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 5238 15206 5290 15258
rect 10918 15206 10970 15258
rect 10982 15206 11034 15258
rect 11046 15206 11098 15258
rect 11110 15206 11162 15258
rect 11174 15206 11226 15258
rect 11238 15206 11290 15258
rect 664 15104 716 15156
rect 1860 15147 1912 15156
rect 1860 15113 1869 15147
rect 1869 15113 1903 15147
rect 1903 15113 1912 15147
rect 1860 15104 1912 15113
rect 2872 15104 2924 15156
rect 3976 15104 4028 15156
rect 5356 15104 5408 15156
rect 6184 15104 6236 15156
rect 7380 15147 7432 15156
rect 7380 15113 7389 15147
rect 7389 15113 7423 15147
rect 7423 15113 7432 15147
rect 7380 15104 7432 15113
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 9496 15104 9548 15156
rect 11704 15104 11756 15156
rect 12808 15104 12860 15156
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 3608 15036 3660 15088
rect 4712 15036 4764 15088
rect 3424 14968 3476 15020
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 4344 14968 4396 15020
rect 3240 14900 3292 14952
rect 6644 14900 6696 14952
rect 7840 14900 7892 14952
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 5448 14832 5500 14884
rect 10692 14764 10744 14816
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 12900 14764 12952 14816
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 13918 14662 13970 14714
rect 13982 14662 14034 14714
rect 14046 14662 14098 14714
rect 14110 14662 14162 14714
rect 14174 14662 14226 14714
rect 14238 14662 14290 14714
rect 1584 14560 1636 14612
rect 8944 14560 8996 14612
rect 9220 14560 9272 14612
rect 3240 14535 3292 14544
rect 3240 14501 3249 14535
rect 3249 14501 3283 14535
rect 3283 14501 3292 14535
rect 3240 14492 3292 14501
rect 1492 14356 1544 14408
rect 3516 14356 3568 14408
rect 8760 14399 8812 14408
rect 8760 14365 8769 14399
rect 8769 14365 8803 14399
rect 8803 14365 8812 14399
rect 8760 14356 8812 14365
rect 2228 14288 2280 14340
rect 5632 14288 5684 14340
rect 8484 14331 8536 14340
rect 8484 14297 8502 14331
rect 8502 14297 8536 14331
rect 8484 14288 8536 14297
rect 4804 14220 4856 14272
rect 6644 14220 6696 14272
rect 9404 14288 9456 14340
rect 10692 14288 10744 14340
rect 11428 14356 11480 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12716 14356 12768 14408
rect 13728 14560 13780 14612
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 11796 14220 11848 14272
rect 12072 14220 12124 14272
rect 12164 14220 12216 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 12624 14220 12676 14272
rect 12900 14220 12952 14272
rect 4918 14118 4970 14170
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 5238 14118 5290 14170
rect 10918 14118 10970 14170
rect 10982 14118 11034 14170
rect 11046 14118 11098 14170
rect 11110 14118 11162 14170
rect 11174 14118 11226 14170
rect 11238 14118 11290 14170
rect 2228 14059 2280 14068
rect 2228 14025 2237 14059
rect 2237 14025 2271 14059
rect 2271 14025 2280 14059
rect 2228 14016 2280 14025
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 2504 13880 2556 13932
rect 2872 13880 2924 13932
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3700 13948 3752 14000
rect 4712 14016 4764 14068
rect 5264 14016 5316 14068
rect 7840 14016 7892 14068
rect 8484 14016 8536 14068
rect 10508 14059 10560 14068
rect 10508 14025 10517 14059
rect 10517 14025 10551 14059
rect 10551 14025 10560 14059
rect 10508 14016 10560 14025
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 11796 14016 11848 14068
rect 12164 14016 12216 14068
rect 1492 13812 1544 13864
rect 3516 13812 3568 13864
rect 4160 13880 4212 13932
rect 4804 13880 4856 13932
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5448 13880 5500 13932
rect 2964 13744 3016 13796
rect 3148 13676 3200 13728
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 4988 13744 5040 13796
rect 5816 13880 5868 13932
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 9864 13948 9916 14000
rect 12624 14016 12676 14068
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 9220 13880 9272 13932
rect 9956 13880 10008 13932
rect 11336 13880 11388 13932
rect 11796 13880 11848 13932
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 9404 13855 9456 13864
rect 9404 13821 9413 13855
rect 9413 13821 9447 13855
rect 9447 13821 9456 13855
rect 9404 13812 9456 13821
rect 10140 13812 10192 13864
rect 11428 13812 11480 13864
rect 11704 13744 11756 13796
rect 3884 13676 3936 13728
rect 3976 13676 4028 13728
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 5172 13676 5224 13728
rect 5632 13676 5684 13728
rect 6552 13676 6604 13728
rect 12440 13812 12492 13864
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 12900 13676 12952 13728
rect 13820 13676 13872 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 13918 13574 13970 13626
rect 13982 13574 14034 13626
rect 14046 13574 14098 13626
rect 14110 13574 14162 13626
rect 14174 13574 14226 13626
rect 14238 13574 14290 13626
rect 3148 13515 3200 13524
rect 3148 13481 3157 13515
rect 3157 13481 3191 13515
rect 3191 13481 3200 13515
rect 3148 13472 3200 13481
rect 3332 13472 3384 13524
rect 5080 13472 5132 13524
rect 5448 13472 5500 13524
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 7840 13472 7892 13524
rect 9680 13472 9732 13524
rect 11428 13472 11480 13524
rect 11704 13472 11756 13524
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 2504 13404 2556 13456
rect 1492 13268 1544 13320
rect 1676 13243 1728 13252
rect 1676 13209 1710 13243
rect 1710 13209 1728 13243
rect 1676 13200 1728 13209
rect 4344 13336 4396 13388
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 3884 13268 3936 13320
rect 3240 13200 3292 13252
rect 3332 13200 3384 13252
rect 3700 13200 3752 13252
rect 4528 13268 4580 13320
rect 2872 13132 2924 13184
rect 2964 13175 3016 13184
rect 2964 13141 2973 13175
rect 2973 13141 3007 13175
rect 3007 13141 3016 13175
rect 2964 13132 3016 13141
rect 4988 13336 5040 13388
rect 6184 13336 6236 13388
rect 6368 13268 6420 13320
rect 8760 13379 8812 13388
rect 8760 13345 8769 13379
rect 8769 13345 8803 13379
rect 8803 13345 8812 13379
rect 8760 13336 8812 13345
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 9772 13268 9824 13320
rect 11336 13268 11388 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 13820 13268 13872 13320
rect 5356 13200 5408 13252
rect 9404 13200 9456 13252
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 5448 13132 5500 13184
rect 7472 13132 7524 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 4918 13030 4970 13082
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 5238 13030 5290 13082
rect 10918 13030 10970 13082
rect 10982 13030 11034 13082
rect 11046 13030 11098 13082
rect 11110 13030 11162 13082
rect 11174 13030 11226 13082
rect 11238 13030 11290 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 5356 12928 5408 12980
rect 6184 12928 6236 12980
rect 4896 12903 4948 12912
rect 4896 12869 4905 12903
rect 4905 12869 4939 12903
rect 4939 12869 4948 12903
rect 4896 12860 4948 12869
rect 1676 12792 1728 12844
rect 6736 12903 6788 12912
rect 6736 12869 6745 12903
rect 6745 12869 6779 12903
rect 6779 12869 6788 12903
rect 6736 12860 6788 12869
rect 8852 12792 8904 12844
rect 9496 12928 9548 12980
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 9128 12792 9180 12844
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 4528 12699 4580 12708
rect 4528 12665 4537 12699
rect 4537 12665 4571 12699
rect 4571 12665 4580 12699
rect 4528 12656 4580 12665
rect 5632 12656 5684 12708
rect 4620 12588 4672 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 11428 12792 11480 12844
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 12440 12928 12492 12980
rect 13820 12928 13872 12980
rect 11980 12792 12032 12844
rect 11796 12656 11848 12708
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 11612 12631 11664 12640
rect 11612 12597 11621 12631
rect 11621 12597 11655 12631
rect 11655 12597 11664 12631
rect 11612 12588 11664 12597
rect 12072 12588 12124 12640
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 13918 12486 13970 12538
rect 13982 12486 14034 12538
rect 14046 12486 14098 12538
rect 14110 12486 14162 12538
rect 14174 12486 14226 12538
rect 14238 12486 14290 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 2872 12384 2924 12436
rect 3516 12384 3568 12436
rect 2320 12248 2372 12300
rect 3056 12248 3108 12300
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3516 12180 3568 12232
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 4436 12316 4488 12368
rect 4712 12316 4764 12368
rect 7104 12384 7156 12436
rect 7748 12384 7800 12436
rect 9220 12384 9272 12436
rect 10692 12384 10744 12436
rect 6736 12248 6788 12300
rect 7840 12248 7892 12300
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 5540 12044 5592 12096
rect 5632 12087 5684 12096
rect 5632 12053 5641 12087
rect 5641 12053 5675 12087
rect 5675 12053 5684 12087
rect 5632 12044 5684 12053
rect 5724 12044 5776 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 7472 12180 7524 12232
rect 7656 12180 7708 12232
rect 10048 12316 10100 12368
rect 10692 12248 10744 12300
rect 7840 12155 7892 12164
rect 7840 12121 7849 12155
rect 7849 12121 7883 12155
rect 7883 12121 7892 12155
rect 7840 12112 7892 12121
rect 8576 12180 8628 12232
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 8852 12180 8904 12232
rect 10232 12180 10284 12232
rect 10416 12223 10468 12232
rect 10416 12189 10426 12223
rect 10426 12189 10460 12223
rect 10460 12189 10468 12223
rect 12164 12384 12216 12436
rect 13084 12384 13136 12436
rect 11520 12316 11572 12368
rect 11612 12248 11664 12300
rect 10416 12180 10468 12189
rect 9312 12112 9364 12164
rect 9588 12155 9640 12164
rect 9588 12121 9597 12155
rect 9597 12121 9631 12155
rect 9631 12121 9640 12155
rect 9588 12112 9640 12121
rect 8024 12044 8076 12096
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 10692 12155 10744 12164
rect 10692 12121 10701 12155
rect 10701 12121 10735 12155
rect 10735 12121 10744 12155
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 10692 12112 10744 12121
rect 11704 12180 11756 12232
rect 12532 12316 12584 12368
rect 13176 12316 13228 12368
rect 13820 12248 13872 12300
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 11796 12044 11848 12096
rect 4918 11942 4970 11994
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 5238 11942 5290 11994
rect 10918 11942 10970 11994
rect 10982 11942 11034 11994
rect 11046 11942 11098 11994
rect 11110 11942 11162 11994
rect 11174 11942 11226 11994
rect 11238 11942 11290 11994
rect 3332 11840 3384 11892
rect 5448 11840 5500 11892
rect 5724 11840 5776 11892
rect 7104 11840 7156 11892
rect 7288 11840 7340 11892
rect 8024 11840 8076 11892
rect 9588 11840 9640 11892
rect 11428 11840 11480 11892
rect 4896 11815 4948 11824
rect 4896 11781 4905 11815
rect 4905 11781 4939 11815
rect 4939 11781 4948 11815
rect 4896 11772 4948 11781
rect 5264 11772 5316 11824
rect 5816 11815 5868 11824
rect 5816 11781 5825 11815
rect 5825 11781 5859 11815
rect 5859 11781 5868 11815
rect 5816 11772 5868 11781
rect 11796 11772 11848 11824
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4436 11704 4488 11756
rect 8484 11704 8536 11756
rect 9128 11704 9180 11756
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 12072 11840 12124 11892
rect 12256 11747 12308 11756
rect 12256 11713 12265 11747
rect 12265 11713 12299 11747
rect 12299 11713 12308 11747
rect 12256 11704 12308 11713
rect 11336 11636 11388 11688
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 12992 11772 13044 11824
rect 13820 11704 13872 11756
rect 10508 11568 10560 11620
rect 12164 11568 12216 11620
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4344 11500 4396 11552
rect 4620 11500 4672 11552
rect 4804 11500 4856 11552
rect 5540 11500 5592 11552
rect 5908 11500 5960 11552
rect 8944 11500 8996 11552
rect 10416 11500 10468 11552
rect 12900 11636 12952 11688
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 13918 11398 13970 11450
rect 13982 11398 14034 11450
rect 14046 11398 14098 11450
rect 14110 11398 14162 11450
rect 14174 11398 14226 11450
rect 14238 11398 14290 11450
rect 3148 11296 3200 11348
rect 4160 11296 4212 11348
rect 5816 11296 5868 11348
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2872 11160 2924 11212
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 2964 11092 3016 11144
rect 3608 11092 3660 11144
rect 3792 11092 3844 11144
rect 4896 11228 4948 11280
rect 4804 11160 4856 11212
rect 4344 11024 4396 11076
rect 2688 10956 2740 11008
rect 3976 10956 4028 11008
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 6736 11228 6788 11280
rect 7564 11228 7616 11280
rect 7748 11271 7800 11280
rect 7748 11237 7757 11271
rect 7757 11237 7791 11271
rect 7791 11237 7800 11271
rect 7748 11228 7800 11237
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 10232 11296 10284 11348
rect 12992 11296 13044 11348
rect 9220 11228 9272 11280
rect 9864 11228 9916 11280
rect 10140 11228 10192 11280
rect 4804 11024 4856 11076
rect 5448 11092 5500 11144
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 6920 11160 6972 11212
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 4620 10999 4672 11008
rect 4620 10965 4629 10999
rect 4629 10965 4663 10999
rect 4663 10965 4672 10999
rect 4620 10956 4672 10965
rect 5264 10956 5316 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 6920 11024 6972 11076
rect 7104 11092 7156 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 7656 11024 7708 11076
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8944 11160 8996 11212
rect 9496 11160 9548 11212
rect 9128 11092 9180 11144
rect 11336 11160 11388 11212
rect 11704 11160 11756 11212
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10140 11092 10192 11144
rect 8760 11067 8812 11076
rect 8760 11033 8769 11067
rect 8769 11033 8803 11067
rect 8803 11033 8812 11067
rect 8760 11024 8812 11033
rect 10784 11067 10836 11076
rect 10784 11033 10793 11067
rect 10793 11033 10827 11067
rect 10827 11033 10836 11067
rect 10784 11024 10836 11033
rect 11060 11092 11112 11144
rect 11796 11092 11848 11144
rect 5724 10956 5776 11008
rect 6460 10956 6512 11008
rect 6736 10956 6788 11008
rect 9036 10956 9088 11008
rect 10692 10956 10744 11008
rect 11888 10956 11940 11008
rect 12532 10956 12584 11008
rect 12716 10956 12768 11008
rect 4918 10854 4970 10906
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 5238 10854 5290 10906
rect 10918 10854 10970 10906
rect 10982 10854 11034 10906
rect 11046 10854 11098 10906
rect 11110 10854 11162 10906
rect 11174 10854 11226 10906
rect 11238 10854 11290 10906
rect 2228 10752 2280 10804
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 2780 10752 2832 10804
rect 3884 10752 3936 10804
rect 4620 10752 4672 10804
rect 5448 10752 5500 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 7932 10752 7984 10804
rect 8668 10752 8720 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 9864 10752 9916 10804
rect 10692 10752 10744 10804
rect 10876 10752 10928 10804
rect 11152 10795 11204 10804
rect 11152 10761 11177 10795
rect 11177 10761 11204 10795
rect 11152 10752 11204 10761
rect 11612 10752 11664 10804
rect 13820 10752 13872 10804
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2596 10616 2648 10668
rect 2504 10548 2556 10600
rect 5632 10684 5684 10736
rect 5908 10684 5960 10736
rect 2872 10616 2924 10668
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4804 10616 4856 10668
rect 6000 10616 6052 10668
rect 6552 10616 6604 10668
rect 3056 10548 3108 10600
rect 4344 10548 4396 10600
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 7104 10616 7156 10668
rect 7288 10616 7340 10668
rect 8484 10616 8536 10668
rect 8576 10616 8628 10668
rect 7196 10548 7248 10600
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9404 10548 9456 10600
rect 5448 10480 5500 10532
rect 9128 10480 9180 10532
rect 10140 10616 10192 10668
rect 10968 10727 11020 10736
rect 10968 10693 10977 10727
rect 10977 10693 11011 10727
rect 11011 10693 11020 10727
rect 10968 10684 11020 10693
rect 11520 10684 11572 10736
rect 11428 10616 11480 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11796 10616 11848 10668
rect 13084 10684 13136 10736
rect 12256 10616 12308 10668
rect 13728 10616 13780 10668
rect 4252 10412 4304 10464
rect 7012 10412 7064 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10876 10412 10928 10464
rect 11060 10412 11112 10464
rect 12532 10591 12584 10600
rect 12532 10557 12541 10591
rect 12541 10557 12575 10591
rect 12575 10557 12584 10591
rect 12532 10548 12584 10557
rect 12808 10412 12860 10464
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 13918 10310 13970 10362
rect 13982 10310 14034 10362
rect 14046 10310 14098 10362
rect 14110 10310 14162 10362
rect 14174 10310 14226 10362
rect 14238 10310 14290 10362
rect 4804 10208 4856 10260
rect 6552 10208 6604 10260
rect 9220 10208 9272 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 2964 10140 3016 10192
rect 1492 10004 1544 10056
rect 7012 10140 7064 10192
rect 8576 10140 8628 10192
rect 11152 10140 11204 10192
rect 6644 10072 6696 10124
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4344 10004 4396 10056
rect 6460 10004 6512 10056
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 1768 9936 1820 9988
rect 3884 9936 3936 9988
rect 3332 9868 3384 9920
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 7840 10072 7892 10124
rect 8944 10072 8996 10124
rect 8576 10004 8628 10056
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 11336 10072 11388 10124
rect 8116 9936 8168 9988
rect 8392 9936 8444 9988
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 12440 9936 12492 9988
rect 13176 9979 13228 9988
rect 13176 9945 13185 9979
rect 13185 9945 13219 9979
rect 13219 9945 13228 9979
rect 13176 9936 13228 9945
rect 13360 9979 13412 9988
rect 13360 9945 13369 9979
rect 13369 9945 13403 9979
rect 13403 9945 13412 9979
rect 13360 9936 13412 9945
rect 13636 9936 13688 9988
rect 6828 9868 6880 9920
rect 8208 9868 8260 9920
rect 9496 9868 9548 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11428 9868 11480 9920
rect 11520 9868 11572 9920
rect 12256 9911 12308 9920
rect 12256 9877 12265 9911
rect 12265 9877 12299 9911
rect 12299 9877 12308 9911
rect 12256 9868 12308 9877
rect 4918 9766 4970 9818
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 5238 9766 5290 9818
rect 10918 9766 10970 9818
rect 10982 9766 11034 9818
rect 11046 9766 11098 9818
rect 11110 9766 11162 9818
rect 11174 9766 11226 9818
rect 11238 9766 11290 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 4252 9664 4304 9716
rect 5448 9664 5500 9716
rect 5540 9664 5592 9716
rect 1860 9596 1912 9648
rect 3056 9528 3108 9580
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 3884 9460 3936 9512
rect 4620 9596 4672 9648
rect 4804 9596 4856 9648
rect 4344 9528 4396 9580
rect 5632 9528 5684 9580
rect 5724 9571 5776 9580
rect 5724 9537 5762 9571
rect 5762 9537 5776 9571
rect 5724 9528 5776 9537
rect 6000 9528 6052 9580
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 6920 9639 6972 9648
rect 6920 9605 6929 9639
rect 6929 9605 6963 9639
rect 6963 9605 6972 9639
rect 6920 9596 6972 9605
rect 7380 9707 7432 9716
rect 7380 9673 7389 9707
rect 7389 9673 7423 9707
rect 7423 9673 7432 9707
rect 7380 9664 7432 9673
rect 7840 9664 7892 9716
rect 10784 9664 10836 9716
rect 12164 9664 12216 9716
rect 12256 9664 12308 9716
rect 12348 9664 12400 9716
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 7196 9528 7248 9580
rect 8116 9596 8168 9648
rect 9404 9596 9456 9648
rect 2504 9392 2556 9444
rect 2872 9392 2924 9444
rect 4068 9392 4120 9444
rect 4804 9392 4856 9444
rect 5356 9392 5408 9444
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 6092 9324 6144 9376
rect 6184 9324 6236 9376
rect 8852 9460 8904 9512
rect 9496 9460 9548 9512
rect 10692 9528 10744 9580
rect 11336 9528 11388 9580
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11888 9528 11940 9580
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 12532 9460 12584 9512
rect 6552 9324 6604 9376
rect 8392 9324 8444 9376
rect 8484 9324 8536 9376
rect 8760 9324 8812 9376
rect 9956 9324 10008 9376
rect 13176 9324 13228 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 13918 9222 13970 9274
rect 13982 9222 14034 9274
rect 14046 9222 14098 9274
rect 14110 9222 14162 9274
rect 14174 9222 14226 9274
rect 14238 9222 14290 9274
rect 2964 9120 3016 9172
rect 3148 9120 3200 9172
rect 4344 9120 4396 9172
rect 5448 9120 5500 9172
rect 6920 9120 6972 9172
rect 8208 9120 8260 9172
rect 9128 9120 9180 9172
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 3056 8984 3108 9036
rect 7196 9052 7248 9104
rect 2688 8916 2740 8968
rect 2964 8916 3016 8968
rect 4620 8984 4672 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 6368 8916 6420 8968
rect 5816 8848 5868 8900
rect 6092 8848 6144 8900
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 3056 8823 3108 8832
rect 3056 8789 3065 8823
rect 3065 8789 3099 8823
rect 3099 8789 3108 8823
rect 3056 8780 3108 8789
rect 6920 8780 6972 8832
rect 7288 8780 7340 8832
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8392 8891 8444 8900
rect 8392 8857 8401 8891
rect 8401 8857 8435 8891
rect 8435 8857 8444 8891
rect 8392 8848 8444 8857
rect 8484 8891 8536 8900
rect 8484 8857 8493 8891
rect 8493 8857 8527 8891
rect 8527 8857 8536 8891
rect 8484 8848 8536 8857
rect 8668 8780 8720 8832
rect 9588 9052 9640 9104
rect 9680 8984 9732 9036
rect 12808 9120 12860 9172
rect 9496 8916 9548 8968
rect 9956 8916 10008 8968
rect 10600 8916 10652 8968
rect 10692 8916 10744 8968
rect 11428 9052 11480 9104
rect 12164 9052 12216 9104
rect 9956 8780 10008 8832
rect 12532 8916 12584 8968
rect 13360 9052 13412 9104
rect 12624 8848 12676 8900
rect 12348 8780 12400 8832
rect 4918 8678 4970 8730
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 5238 8678 5290 8730
rect 10918 8678 10970 8730
rect 10982 8678 11034 8730
rect 11046 8678 11098 8730
rect 11110 8678 11162 8730
rect 11174 8678 11226 8730
rect 11238 8678 11290 8730
rect 2504 8576 2556 8628
rect 3056 8576 3108 8628
rect 3332 8576 3384 8628
rect 4804 8576 4856 8628
rect 6000 8576 6052 8628
rect 2964 8508 3016 8560
rect 4344 8508 4396 8560
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 6736 8508 6788 8560
rect 9772 8576 9824 8628
rect 6184 8372 6236 8424
rect 7288 8440 7340 8492
rect 8392 8440 8444 8492
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 6828 8372 6880 8424
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 12256 8576 12308 8628
rect 10140 8508 10192 8560
rect 11704 8508 11756 8560
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 13360 8508 13412 8560
rect 11060 8372 11112 8424
rect 11612 8372 11664 8424
rect 11336 8304 11388 8356
rect 2320 8279 2372 8288
rect 2320 8245 2329 8279
rect 2329 8245 2363 8279
rect 2363 8245 2372 8279
rect 2320 8236 2372 8245
rect 5448 8279 5500 8288
rect 5448 8245 5457 8279
rect 5457 8245 5491 8279
rect 5491 8245 5500 8279
rect 5448 8236 5500 8245
rect 6092 8236 6144 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 9036 8236 9088 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 13918 8134 13970 8186
rect 13982 8134 14034 8186
rect 14046 8134 14098 8186
rect 14110 8134 14162 8186
rect 14174 8134 14226 8186
rect 14238 8134 14290 8186
rect 4160 8075 4212 8084
rect 4160 8041 4169 8075
rect 4169 8041 4203 8075
rect 4203 8041 4212 8075
rect 4160 8032 4212 8041
rect 4528 8032 4580 8084
rect 1492 7896 1544 7948
rect 2596 7828 2648 7880
rect 3332 7828 3384 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4712 7828 4764 7880
rect 6000 8032 6052 8084
rect 6552 8032 6604 8084
rect 7380 8032 7432 8084
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 9864 8032 9916 8084
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 5540 7964 5592 8016
rect 6184 7964 6236 8016
rect 5448 7896 5500 7948
rect 9404 7964 9456 8016
rect 10232 7964 10284 8016
rect 11060 8007 11112 8016
rect 11060 7973 11069 8007
rect 11069 7973 11103 8007
rect 11103 7973 11112 8007
rect 11060 7964 11112 7973
rect 6920 7896 6972 7948
rect 7196 7896 7248 7948
rect 7288 7896 7340 7948
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 2320 7803 2372 7812
rect 2320 7769 2354 7803
rect 2354 7769 2372 7803
rect 2320 7760 2372 7769
rect 3884 7692 3936 7744
rect 4068 7692 4120 7744
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 7012 7828 7064 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8484 7828 8536 7880
rect 9036 7828 9088 7880
rect 9680 7828 9732 7880
rect 5632 7692 5684 7744
rect 7840 7692 7892 7744
rect 8392 7692 8444 7744
rect 9588 7760 9640 7812
rect 10692 7828 10744 7880
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 11888 7828 11940 7880
rect 10140 7692 10192 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 4918 7590 4970 7642
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 5238 7590 5290 7642
rect 10918 7590 10970 7642
rect 10982 7590 11034 7642
rect 11046 7590 11098 7642
rect 11110 7590 11162 7642
rect 11174 7590 11226 7642
rect 11238 7590 11290 7642
rect 3332 7488 3384 7540
rect 4160 7488 4212 7540
rect 5540 7488 5592 7540
rect 3792 7420 3844 7472
rect 3424 7352 3476 7404
rect 7012 7488 7064 7540
rect 6092 7463 6144 7472
rect 6092 7429 6101 7463
rect 6101 7429 6135 7463
rect 6135 7429 6144 7463
rect 6092 7420 6144 7429
rect 7104 7420 7156 7472
rect 10508 7488 10560 7540
rect 6000 7352 6052 7404
rect 6460 7352 6512 7404
rect 6736 7352 6788 7404
rect 5816 7284 5868 7336
rect 7748 7284 7800 7336
rect 9496 7420 9548 7472
rect 9956 7420 10008 7472
rect 10232 7420 10284 7472
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 3884 7216 3936 7268
rect 6460 7216 6512 7268
rect 9312 7284 9364 7336
rect 9496 7284 9548 7336
rect 11336 7420 11388 7472
rect 10692 7216 10744 7268
rect 4068 7148 4120 7200
rect 5724 7148 5776 7200
rect 7472 7148 7524 7200
rect 7840 7148 7892 7200
rect 8576 7148 8628 7200
rect 10048 7148 10100 7200
rect 10140 7148 10192 7200
rect 11060 7148 11112 7200
rect 11796 7148 11848 7200
rect 12624 7148 12676 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 13918 7046 13970 7098
rect 13982 7046 14034 7098
rect 14046 7046 14098 7098
rect 14110 7046 14162 7098
rect 14174 7046 14226 7098
rect 14238 7046 14290 7098
rect 3424 6944 3476 6996
rect 4712 6944 4764 6996
rect 7840 6944 7892 6996
rect 8392 6944 8444 6996
rect 9588 6944 9640 6996
rect 9864 6944 9916 6996
rect 10324 6944 10376 6996
rect 11060 6944 11112 6996
rect 4804 6876 4856 6928
rect 2596 6808 2648 6860
rect 4344 6740 4396 6792
rect 4252 6672 4304 6724
rect 7196 6876 7248 6928
rect 9496 6876 9548 6928
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 5632 6672 5684 6724
rect 7472 6740 7524 6792
rect 8024 6740 8076 6792
rect 6368 6672 6420 6724
rect 5448 6604 5500 6656
rect 5816 6604 5868 6656
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 10232 6740 10284 6792
rect 10692 6740 10744 6792
rect 11888 6944 11940 6996
rect 12256 6944 12308 6996
rect 9772 6604 9824 6656
rect 10784 6604 10836 6656
rect 12624 6740 12676 6792
rect 11336 6672 11388 6724
rect 12164 6604 12216 6656
rect 12256 6604 12308 6656
rect 4918 6502 4970 6554
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 5238 6502 5290 6554
rect 10918 6502 10970 6554
rect 10982 6502 11034 6554
rect 11046 6502 11098 6554
rect 11110 6502 11162 6554
rect 11174 6502 11226 6554
rect 11238 6502 11290 6554
rect 8484 6443 8536 6452
rect 8484 6409 8493 6443
rect 8493 6409 8527 6443
rect 8527 6409 8536 6443
rect 8484 6400 8536 6409
rect 2412 6332 2464 6384
rect 7748 6332 7800 6384
rect 8024 6375 8076 6384
rect 8024 6341 8033 6375
rect 8033 6341 8067 6375
rect 8067 6341 8076 6375
rect 8024 6332 8076 6341
rect 9864 6332 9916 6384
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 1676 6196 1728 6248
rect 4068 6196 4120 6248
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 5448 6196 5500 6248
rect 1584 6060 1636 6112
rect 4252 6128 4304 6180
rect 8392 6264 8444 6316
rect 8576 6264 8628 6316
rect 10232 6400 10284 6452
rect 11336 6400 11388 6452
rect 9772 6171 9824 6180
rect 9772 6137 9781 6171
rect 9781 6137 9815 6171
rect 9815 6137 9824 6171
rect 9772 6128 9824 6137
rect 10692 6264 10744 6316
rect 10048 6196 10100 6248
rect 10324 6239 10376 6248
rect 10324 6205 10333 6239
rect 10333 6205 10367 6239
rect 10367 6205 10376 6239
rect 10324 6196 10376 6205
rect 10232 6128 10284 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 6092 6060 6144 6112
rect 7840 6060 7892 6112
rect 9588 6060 9640 6112
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11704 6196 11756 6248
rect 10876 6128 10928 6180
rect 12072 6239 12124 6248
rect 12072 6205 12081 6239
rect 12081 6205 12115 6239
rect 12115 6205 12124 6239
rect 12072 6196 12124 6205
rect 13820 6400 13872 6452
rect 12624 6332 12676 6384
rect 12348 6196 12400 6248
rect 12808 6196 12860 6248
rect 14464 6196 14516 6248
rect 11612 6060 11664 6112
rect 12900 6128 12952 6180
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 13918 5958 13970 6010
rect 13982 5958 14034 6010
rect 14046 5958 14098 6010
rect 14110 5958 14162 6010
rect 14174 5958 14226 6010
rect 14238 5958 14290 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 3424 5856 3476 5908
rect 3608 5856 3660 5908
rect 5540 5856 5592 5908
rect 5908 5856 5960 5908
rect 8392 5856 8444 5908
rect 6276 5788 6328 5840
rect 5172 5720 5224 5772
rect 3608 5584 3660 5636
rect 4252 5652 4304 5704
rect 4528 5652 4580 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 5632 5584 5684 5636
rect 5816 5516 5868 5568
rect 6552 5584 6604 5636
rect 8484 5788 8536 5840
rect 9220 5856 9272 5908
rect 9404 5856 9456 5908
rect 10876 5856 10928 5908
rect 11152 5856 11204 5908
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 11796 5856 11848 5908
rect 12072 5856 12124 5908
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 9588 5788 9640 5840
rect 10232 5788 10284 5840
rect 10600 5788 10652 5840
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 7840 5627 7892 5636
rect 7104 5516 7156 5568
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 9772 5652 9824 5704
rect 10048 5720 10100 5772
rect 10140 5763 10192 5772
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 10784 5652 10836 5704
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 12072 5720 12124 5772
rect 10508 5584 10560 5636
rect 10600 5584 10652 5636
rect 10968 5584 11020 5636
rect 12348 5652 12400 5704
rect 12624 5652 12676 5704
rect 12808 5695 12860 5704
rect 12808 5661 12842 5695
rect 12842 5661 12860 5695
rect 12808 5652 12860 5661
rect 11888 5627 11940 5636
rect 11888 5593 11897 5627
rect 11897 5593 11931 5627
rect 11931 5593 11940 5627
rect 11888 5584 11940 5593
rect 11980 5584 12032 5636
rect 13544 5584 13596 5636
rect 10784 5516 10836 5568
rect 11428 5516 11480 5568
rect 13820 5516 13872 5568
rect 14556 5516 14608 5568
rect 4918 5414 4970 5466
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 5238 5414 5290 5466
rect 10918 5414 10970 5466
rect 10982 5414 11034 5466
rect 11046 5414 11098 5466
rect 11110 5414 11162 5466
rect 11174 5414 11226 5466
rect 11238 5414 11290 5466
rect 2320 5176 2372 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4528 5312 4580 5364
rect 8760 5312 8812 5364
rect 9312 5312 9364 5364
rect 9496 5312 9548 5364
rect 11796 5312 11848 5364
rect 6092 5244 6144 5296
rect 4436 5176 4488 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 8300 5244 8352 5296
rect 10416 5244 10468 5296
rect 6736 5176 6788 5185
rect 4160 5040 4212 5092
rect 3332 4972 3384 5024
rect 4068 4972 4120 5024
rect 5816 4972 5868 5024
rect 6828 5108 6880 5160
rect 9588 5176 9640 5228
rect 10784 5176 10836 5228
rect 10968 5176 11020 5228
rect 12716 5312 12768 5364
rect 12900 5312 12952 5364
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 12348 5176 12400 5228
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 12716 5108 12768 5117
rect 6644 4972 6696 5024
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 8392 4972 8444 5024
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 10968 4972 11020 5024
rect 12256 4972 12308 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 13918 4870 13970 4922
rect 13982 4870 14034 4922
rect 14046 4870 14098 4922
rect 14110 4870 14162 4922
rect 14174 4870 14226 4922
rect 14238 4870 14290 4922
rect 8852 4768 8904 4820
rect 10784 4768 10836 4820
rect 11888 4768 11940 4820
rect 9312 4700 9364 4752
rect 3700 4632 3752 4684
rect 1676 4564 1728 4616
rect 2044 4496 2096 4548
rect 2320 4428 2372 4480
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 8484 4564 8536 4616
rect 8576 4564 8628 4616
rect 9220 4607 9272 4616
rect 4160 4539 4212 4548
rect 4160 4505 4169 4539
rect 4169 4505 4203 4539
rect 4203 4505 4212 4539
rect 4160 4496 4212 4505
rect 4804 4496 4856 4548
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 8944 4539 8996 4548
rect 8944 4505 8953 4539
rect 8953 4505 8987 4539
rect 8987 4505 8996 4539
rect 8944 4496 8996 4505
rect 12624 4564 12676 4616
rect 10508 4496 10560 4548
rect 10784 4496 10836 4548
rect 12256 4539 12308 4548
rect 12256 4505 12297 4539
rect 12297 4505 12308 4539
rect 12256 4496 12308 4505
rect 12808 4539 12860 4548
rect 12808 4505 12842 4539
rect 12842 4505 12860 4539
rect 12808 4496 12860 4505
rect 4620 4428 4672 4480
rect 6736 4428 6788 4480
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 8300 4428 8352 4480
rect 9404 4428 9456 4480
rect 10324 4428 10376 4480
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 13820 4428 13872 4480
rect 14372 4428 14424 4480
rect 4918 4326 4970 4378
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 5238 4326 5290 4378
rect 10918 4326 10970 4378
rect 10982 4326 11034 4378
rect 11046 4326 11098 4378
rect 11110 4326 11162 4378
rect 11174 4326 11226 4378
rect 11238 4326 11290 4378
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 3792 4224 3844 4276
rect 3976 4224 4028 4276
rect 3332 4088 3384 4140
rect 4804 4156 4856 4208
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4068 4020 4120 4072
rect 3148 3952 3200 4004
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 6828 4224 6880 4276
rect 7012 4224 7064 4276
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 9312 4224 9364 4276
rect 9772 4224 9824 4276
rect 12440 4224 12492 4276
rect 12808 4267 12860 4276
rect 12808 4233 12817 4267
rect 12817 4233 12851 4267
rect 12851 4233 12860 4267
rect 12808 4224 12860 4233
rect 13176 4224 13228 4276
rect 6736 4199 6788 4208
rect 6736 4165 6745 4199
rect 6745 4165 6779 4199
rect 6779 4165 6788 4199
rect 6736 4156 6788 4165
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 8392 4199 8444 4208
rect 8392 4165 8401 4199
rect 8401 4165 8435 4199
rect 8435 4165 8444 4199
rect 8392 4156 8444 4165
rect 8300 4088 8352 4140
rect 9036 4131 9088 4140
rect 9036 4097 9045 4131
rect 9045 4097 9079 4131
rect 9079 4097 9088 4131
rect 9036 4088 9088 4097
rect 9220 4088 9272 4140
rect 9404 4156 9456 4208
rect 9680 4156 9732 4208
rect 9864 4199 9916 4208
rect 9864 4165 9873 4199
rect 9873 4165 9907 4199
rect 9907 4165 9916 4199
rect 9864 4156 9916 4165
rect 5448 3952 5500 4004
rect 7104 4020 7156 4072
rect 9128 4020 9180 4072
rect 10692 4088 10744 4140
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 9864 4020 9916 4072
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10600 4020 10652 4072
rect 8852 3952 8904 4004
rect 9772 3952 9824 4004
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 7840 3884 7892 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 10048 3884 10100 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 13918 3782 13970 3834
rect 13982 3782 14034 3834
rect 14046 3782 14098 3834
rect 14110 3782 14162 3834
rect 14174 3782 14226 3834
rect 14238 3782 14290 3834
rect 3240 3680 3292 3732
rect 4804 3680 4856 3732
rect 4896 3680 4948 3732
rect 5632 3680 5684 3732
rect 5448 3544 5500 3596
rect 6368 3680 6420 3732
rect 7380 3680 7432 3732
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 5816 3476 5868 3528
rect 8392 3476 8444 3528
rect 9036 3476 9088 3528
rect 10508 3476 10560 3528
rect 6368 3408 6420 3460
rect 10600 3408 10652 3460
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 4160 3340 4212 3392
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 6920 3340 6972 3392
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 4918 3238 4970 3290
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 5238 3238 5290 3290
rect 10918 3238 10970 3290
rect 10982 3238 11034 3290
rect 11046 3238 11098 3290
rect 11110 3238 11162 3290
rect 11174 3238 11226 3290
rect 11238 3238 11290 3290
rect 4252 3136 4304 3188
rect 5632 3136 5684 3188
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 9036 3136 9088 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 14464 3136 14516 3188
rect 1676 3000 1728 3052
rect 3792 3000 3844 3052
rect 5816 3068 5868 3120
rect 7104 3068 7156 3120
rect 4896 3043 4948 3052
rect 4896 3009 4930 3043
rect 4930 3009 4948 3043
rect 4896 3000 4948 3009
rect 5908 3000 5960 3052
rect 7840 3068 7892 3120
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 13452 3000 13504 3052
rect 11060 2796 11112 2848
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 13918 2694 13970 2746
rect 13982 2694 14034 2746
rect 14046 2694 14098 2746
rect 14110 2694 14162 2746
rect 14174 2694 14226 2746
rect 14238 2694 14290 2746
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4252 2592 4304 2644
rect 1676 2456 1728 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2320 2388 2372 2440
rect 2504 2431 2556 2440
rect 2504 2397 2538 2431
rect 2538 2397 2556 2431
rect 2504 2388 2556 2397
rect 4160 2388 4212 2440
rect 4344 2388 4396 2440
rect 4896 2592 4948 2644
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 7104 2456 7156 2508
rect 5632 2388 5684 2440
rect 6000 2388 6052 2440
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7472 2431 7524 2440
rect 7472 2397 7506 2431
rect 7506 2397 7524 2431
rect 7472 2388 7524 2397
rect 8760 2388 8812 2440
rect 10324 2388 10376 2440
rect 10508 2592 10560 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 11060 2456 11112 2508
rect 14372 2456 14424 2508
rect 9312 2320 9364 2372
rect 9772 2320 9824 2372
rect 14464 2388 14516 2440
rect 756 2252 808 2304
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 3700 2252 3752 2304
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 8668 2252 8720 2304
rect 14924 2320 14976 2372
rect 11336 2252 11388 2304
rect 12348 2252 12400 2304
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 4918 2150 4970 2202
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 5238 2150 5290 2202
rect 10918 2150 10970 2202
rect 10982 2150 11034 2202
rect 11046 2150 11098 2202
rect 11110 2150 11162 2202
rect 11174 2150 11226 2202
rect 11238 2150 11290 2202
<< metal2 >>
rect 662 17064 718 17864
rect 1766 17218 1822 17864
rect 1766 17190 1900 17218
rect 1766 17064 1822 17190
rect 676 15162 704 17064
rect 1872 15162 1900 17190
rect 2870 17064 2926 17864
rect 3974 17064 4030 17864
rect 5078 17064 5134 17864
rect 6182 17064 6238 17864
rect 7286 17218 7342 17864
rect 8390 17218 8446 17864
rect 7286 17190 7420 17218
rect 7286 17064 7342 17190
rect 2884 15162 2912 17064
rect 3988 15162 4016 17064
rect 5092 15994 5120 17064
rect 5092 15966 5396 15994
rect 4916 15260 5292 15269
rect 4972 15258 4996 15260
rect 5052 15258 5076 15260
rect 5132 15258 5156 15260
rect 5212 15258 5236 15260
rect 4972 15206 4982 15258
rect 5226 15206 5236 15258
rect 4972 15204 4996 15206
rect 5052 15204 5076 15206
rect 5132 15204 5156 15206
rect 5212 15204 5236 15206
rect 4916 15195 5292 15204
rect 5368 15162 5396 15966
rect 6196 15162 6224 17064
rect 7392 15162 7420 17190
rect 8390 17190 8524 17218
rect 8390 17064 8446 17190
rect 8496 15162 8524 17190
rect 9494 17064 9550 17864
rect 10598 17064 10654 17864
rect 11702 17064 11758 17864
rect 12806 17064 12862 17864
rect 13910 17064 13966 17864
rect 15014 17064 15070 17864
rect 9508 15162 9536 17064
rect 664 15156 716 15162
rect 664 15098 716 15104
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 1596 14618 1624 14962
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 3252 14550 3280 14894
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1504 13870 1532 14350
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 2240 14074 2268 14282
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2226 13968 2282 13977
rect 2504 13932 2556 13938
rect 2282 13912 2360 13920
rect 2226 13903 2228 13912
rect 2280 13892 2360 13912
rect 2228 13874 2280 13880
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13326 1532 13806
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 10062 1532 13262
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 12986 1716 13194
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12442 1716 12786
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 2332 12306 2360 13892
rect 2504 13874 2556 13880
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2516 13462 2544 13874
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10146 1808 11154
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10810 2268 11018
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2332 10674 2360 12242
rect 2516 12238 2544 13398
rect 2884 13326 2912 13874
rect 2976 13802 3004 13874
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2872 13320 2924 13326
rect 3068 13274 3096 13874
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13530 3188 13670
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2872 13262 2924 13268
rect 2976 13246 3096 13274
rect 3252 13258 3280 14486
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 13530 3372 13670
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3240 13252 3292 13258
rect 2976 13190 3004 13246
rect 3240 13194 3292 13200
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2884 12442 2912 13126
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2976 12434 3004 13126
rect 2976 12406 3096 12434
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2516 10606 2544 12174
rect 2976 11370 3004 12406
rect 3068 12306 3096 12406
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2792 11342 3004 11370
rect 3160 11354 3188 12174
rect 3148 11348 3200 11354
rect 2688 11144 2740 11150
rect 2792 11098 2820 11342
rect 3148 11290 3200 11296
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2740 11092 2820 11098
rect 2688 11086 2820 11092
rect 2700 11070 2820 11086
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2700 10810 2728 10950
rect 2792 10810 2820 11070
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2884 10674 2912 11154
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 1780 10118 1900 10146
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 7954 1532 9998
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9722 1808 9930
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1872 9654 1900 10118
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 2516 9450 2544 10542
rect 2608 9674 2636 10610
rect 2976 10198 3004 11086
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2608 9646 2728 9674
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 2700 8974 2728 9646
rect 3068 9586 3096 10542
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9042 2912 9386
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3068 9042 3096 9522
rect 3160 9178 3188 9522
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8634 2544 8774
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2976 8566 3004 8910
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8634 3096 8774
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2320 8288 2372 8294
rect 3252 8276 3280 13194
rect 3344 11898 3372 13194
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9518 3372 9862
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 8634 3372 9454
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2320 8230 2372 8236
rect 3160 8248 3280 8276
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 2332 7818 2360 8230
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2608 6866 2636 7822
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 2446 1624 6054
rect 1688 4622 1716 6190
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 2424 5914 2452 6326
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 3058 1716 4558
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 2056 4282 2084 4490
rect 2332 4486 2360 5170
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 2514 1716 2994
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 2332 2446 2360 4422
rect 3160 4010 3188 8248
rect 3344 7886 3372 8570
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7546 3372 7822
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3436 7410 3464 14962
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3528 13870 3556 14350
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3528 12238 3556 12378
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 7002 3464 7346
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3344 4146 3372 4966
rect 3528 4570 3556 12174
rect 3620 11150 3648 15030
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3712 13818 3740 13942
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3712 13790 4016 13818
rect 3988 13734 4016 13790
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3896 13326 3924 13670
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3620 5914 3648 6258
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3620 5234 3648 5578
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 4690 3740 13194
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10674 3832 11086
rect 3896 10810 3924 13262
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11665 4016 11698
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3884 10668 3936 10674
rect 3988 10656 4016 10950
rect 3936 10628 4016 10656
rect 3884 10610 3936 10616
rect 3896 9994 3924 10610
rect 4080 10062 4108 12038
rect 4172 11642 4200 13874
rect 4264 12434 4292 14962
rect 4356 13394 4384 14962
rect 4724 14074 4752 15030
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 14068 4764 14074
rect 4540 14028 4712 14056
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4540 13326 4568 14028
rect 4712 14010 4764 14016
rect 4816 13938 4844 14214
rect 4916 14172 5292 14181
rect 4972 14170 4996 14172
rect 5052 14170 5076 14172
rect 5132 14170 5156 14172
rect 5212 14170 5236 14172
rect 4972 14118 4982 14170
rect 5226 14118 5236 14170
rect 4972 14116 4996 14118
rect 5052 14116 5076 14118
rect 5132 14116 5156 14118
rect 5212 14116 5236 14118
rect 4916 14107 5292 14116
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5276 13938 5304 14010
rect 5460 13938 5488 14826
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5000 13394 5028 13738
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5092 13530 5120 13670
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 5184 13190 5212 13670
rect 5276 13190 5304 13874
rect 5368 13258 5396 13874
rect 5644 13818 5672 14282
rect 6656 14278 6684 14894
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 7852 14074 7880 14894
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8496 14074 8524 14282
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 5460 13790 5672 13818
rect 5460 13530 5488 13790
rect 5632 13728 5684 13734
rect 5828 13682 5856 13874
rect 5684 13676 5856 13682
rect 5632 13670 5856 13676
rect 5644 13654 5856 13670
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 6196 13394 6224 13874
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6564 13530 6592 13670
rect 7852 13530 7880 14010
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 8772 13394 8800 14350
rect 8956 13938 8984 14554
rect 9232 13977 9260 14554
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9218 13968 9274 13977
rect 8944 13932 8996 13938
rect 9218 13903 9220 13912
rect 8944 13874 8996 13880
rect 9272 13903 9274 13912
rect 9220 13874 9272 13880
rect 9416 13870 9444 14282
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4916 13084 5292 13093
rect 4972 13082 4996 13084
rect 5052 13082 5076 13084
rect 5132 13082 5156 13084
rect 5212 13082 5236 13084
rect 4972 13030 4982 13082
rect 5226 13030 5236 13082
rect 4972 13028 4996 13030
rect 5052 13028 5076 13030
rect 5132 13028 5156 13030
rect 5212 13028 5236 13030
rect 4916 13019 5292 13028
rect 5368 12986 5396 13194
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4264 12406 4476 12434
rect 4448 12374 4476 12406
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4434 11792 4490 11801
rect 4434 11727 4436 11736
rect 4488 11727 4490 11736
rect 4436 11698 4488 11704
rect 4172 11614 4476 11642
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4172 11354 4200 11494
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4356 11082 4384 11494
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 4264 9926 4292 10406
rect 4356 10062 4384 10542
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4264 9722 4292 9862
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4356 9586 4384 9998
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 7478 3832 7822
rect 3896 7750 3924 9454
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4080 7750 4108 9386
rect 4356 9178 4384 9522
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3896 7274 3924 7686
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 4080 7206 4108 7686
rect 4172 7546 4200 8026
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4264 6730 4292 7686
rect 4356 6798 4384 8502
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5030 4108 6190
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4264 5710 4292 6122
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4172 5098 4200 5578
rect 4448 5234 4476 11614
rect 4540 8974 4568 12650
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4632 12102 4660 12582
rect 4908 12434 4936 12854
rect 5460 12434 5488 13126
rect 6196 12986 6224 13330
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 4816 12406 4936 12434
rect 5368 12406 5488 12434
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11558 4660 12038
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4632 10810 4660 10950
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4724 10690 4752 12310
rect 4816 11558 4844 12406
rect 4916 11996 5292 12005
rect 4972 11994 4996 11996
rect 5052 11994 5076 11996
rect 5132 11994 5156 11996
rect 5212 11994 5236 11996
rect 4972 11942 4982 11994
rect 5226 11942 5236 11994
rect 4972 11940 4996 11942
rect 5052 11940 5076 11942
rect 5132 11940 5156 11942
rect 5212 11940 5236 11942
rect 4916 11931 5292 11940
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4908 11286 4936 11766
rect 4896 11280 4948 11286
rect 4896 11222 4948 11228
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 11082 4844 11154
rect 4896 11144 4948 11150
rect 4894 11112 4896 11121
rect 4948 11112 4950 11121
rect 4804 11076 4856 11082
rect 4894 11047 4950 11056
rect 4804 11018 4856 11024
rect 4632 10662 4752 10690
rect 4816 10674 4844 11018
rect 5276 11014 5304 11766
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 4916 10908 5292 10917
rect 4972 10906 4996 10908
rect 5052 10906 5076 10908
rect 5132 10906 5156 10908
rect 5212 10906 5236 10908
rect 4972 10854 4982 10906
rect 5226 10854 5236 10906
rect 4972 10852 4996 10854
rect 5052 10852 5076 10854
rect 5132 10852 5156 10854
rect 5212 10852 5236 10854
rect 4916 10843 5292 10852
rect 4804 10668 4856 10674
rect 4632 9654 4660 10662
rect 4804 10610 4856 10616
rect 4816 10266 4844 10610
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4816 9654 4844 10202
rect 4916 9820 5292 9829
rect 4972 9818 4996 9820
rect 5052 9818 5076 9820
rect 5132 9818 5156 9820
rect 5212 9818 5236 9820
rect 4972 9766 4982 9818
rect 5226 9766 5236 9818
rect 4972 9764 4996 9766
rect 5052 9764 5076 9766
rect 5132 9764 5156 9766
rect 5212 9764 5236 9766
rect 4916 9755 5292 9764
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4632 9042 4660 9454
rect 5368 9450 5396 12406
rect 5644 12102 5672 12650
rect 6380 12434 6408 13262
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6288 12406 6408 12434
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5460 11150 5488 11834
rect 5552 11558 5580 12038
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5460 10810 5488 10950
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5644 10742 5672 12038
rect 5736 11898 5764 12038
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5736 11665 5764 11834
rect 5816 11824 5868 11830
rect 6012 11801 6040 12038
rect 5816 11766 5868 11772
rect 5998 11792 6054 11801
rect 5722 11656 5778 11665
rect 5722 11591 5778 11600
rect 5736 11014 5764 11591
rect 5828 11354 5856 11766
rect 5998 11727 6054 11736
rect 5908 11552 5960 11558
rect 6012 11540 6040 11727
rect 5960 11512 6040 11540
rect 5908 11494 5960 11500
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5920 11234 5948 11494
rect 5828 11206 5948 11234
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 9722 5488 10474
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5540 9716 5592 9722
rect 5828 9674 5856 11206
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5920 10742 5948 11086
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 6012 10674 6040 11086
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5540 9658 5592 9664
rect 5552 9602 5580 9658
rect 5460 9574 5580 9602
rect 5644 9646 5856 9674
rect 5644 9586 5672 9646
rect 5632 9580 5684 9586
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8090 4568 8910
rect 4816 8634 4844 9386
rect 5460 9178 5488 9574
rect 5632 9522 5684 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 4916 8732 5292 8741
rect 4972 8730 4996 8732
rect 5052 8730 5076 8732
rect 5132 8730 5156 8732
rect 5212 8730 5236 8732
rect 4972 8678 4982 8730
rect 5226 8678 5236 8730
rect 4972 8676 4996 8678
rect 5052 8676 5076 8678
rect 5132 8676 5156 8678
rect 5212 8676 5236 8678
rect 4916 8667 5292 8676
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 5460 7954 5488 8230
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 4712 7880 4764 7886
rect 4764 7840 4844 7868
rect 4712 7822 4764 7828
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4724 5710 4752 6938
rect 4816 6934 4844 7840
rect 4916 7644 5292 7653
rect 4972 7642 4996 7644
rect 5052 7642 5076 7644
rect 5132 7642 5156 7644
rect 5212 7642 5236 7644
rect 4972 7590 4982 7642
rect 5226 7590 5236 7642
rect 4972 7588 4996 7590
rect 5052 7588 5076 7590
rect 5132 7588 5156 7590
rect 5212 7588 5236 7590
rect 4916 7579 5292 7588
rect 5552 7546 5580 7958
rect 5644 7750 5672 9522
rect 5736 8498 5764 9522
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5828 8786 5856 8842
rect 6012 8786 6040 9522
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6104 8906 6132 9318
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 5828 8758 6040 8786
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5828 7342 5856 8758
rect 6012 8634 6040 8758
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6196 8430 6224 9318
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6012 7410 6040 8026
rect 6104 7478 6132 8230
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6196 7886 6224 7958
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 5736 6798 5764 7142
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5816 6792 5868 6798
rect 5868 6740 5948 6746
rect 5816 6734 5948 6740
rect 5632 6724 5684 6730
rect 5828 6718 5948 6734
rect 5632 6666 5684 6672
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4916 6556 5292 6565
rect 4972 6554 4996 6556
rect 5052 6554 5076 6556
rect 5132 6554 5156 6556
rect 5212 6554 5236 6556
rect 4972 6502 4982 6554
rect 5226 6502 5236 6554
rect 4972 6500 4996 6502
rect 5052 6500 5076 6502
rect 5132 6500 5156 6502
rect 5212 6500 5236 6502
rect 4916 6491 5292 6500
rect 5460 6254 5488 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5184 5778 5212 6190
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4540 5370 4568 5646
rect 4916 5468 5292 5477
rect 4972 5466 4996 5468
rect 5052 5466 5076 5468
rect 5132 5466 5156 5468
rect 5212 5466 5236 5468
rect 4972 5414 4982 5466
rect 5226 5414 5236 5466
rect 4972 5412 4996 5414
rect 5052 5412 5076 5414
rect 5132 5412 5156 5414
rect 5212 5412 5236 5414
rect 4916 5403 5292 5412
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3528 4542 3924 4570
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4282 3832 4422
rect 3792 4276 3844 4282
rect 3896 4264 3924 4542
rect 3976 4276 4028 4282
rect 3896 4236 3976 4264
rect 3792 4218 3844 4224
rect 3976 4218 4028 4224
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 4080 4078 4108 4966
rect 4172 4554 4200 5034
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3738 3280 3878
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 2700 2774 2728 3334
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 2516 2746 2728 2774
rect 2516 2446 2544 2746
rect 3804 2650 3832 2994
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4172 2446 4200 3334
rect 4264 3194 4292 4082
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4264 2650 4292 3130
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4356 2446 4384 4558
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4146 4660 4422
rect 4816 4214 4844 4490
rect 4916 4380 5292 4389
rect 4972 4378 4996 4380
rect 5052 4378 5076 4380
rect 5132 4378 5156 4380
rect 5212 4378 5236 4380
rect 4972 4326 4982 4378
rect 5226 4326 5236 4378
rect 4972 4324 4996 4326
rect 5052 4324 5076 4326
rect 5132 4324 5156 4326
rect 5212 4324 5236 4326
rect 4916 4315 5292 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3738 4844 3878
rect 4908 3738 4936 4082
rect 5460 4010 5488 6190
rect 5552 5914 5580 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5642 5672 6666
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5828 5574 5856 6598
rect 5920 5914 5948 6718
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5030 5856 5510
rect 6104 5302 6132 6054
rect 6288 5846 6316 12406
rect 6748 12306 6776 12854
rect 7484 12594 7512 13126
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8760 12640 8812 12646
rect 7484 12566 7880 12594
rect 8760 12582 8812 12588
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11286 6776 12242
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6932 11218 6960 12174
rect 7116 11898 7144 12378
rect 7484 12238 7512 12566
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6644 11144 6696 11150
rect 6828 11144 6880 11150
rect 6644 11086 6696 11092
rect 6748 11104 6828 11132
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10810 6500 10950
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6564 10674 6592 11086
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 10266 6592 10610
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6380 7886 6408 8910
rect 6472 7970 6500 9998
rect 6564 9382 6592 10202
rect 6656 10130 6684 11086
rect 6748 11014 6776 11104
rect 6828 11086 6880 11092
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10674 6776 10950
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9586 6684 10066
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6748 8566 6776 10610
rect 6932 10130 6960 11018
rect 7116 10674 7144 11086
rect 7300 10674 7328 11834
rect 7484 11268 7512 12174
rect 7564 11280 7616 11286
rect 7484 11240 7564 11268
rect 7564 11222 7616 11228
rect 7668 11082 7696 12174
rect 7760 11286 7788 12378
rect 7852 12306 7880 12566
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 8772 12434 8800 12582
rect 8680 12406 8800 12434
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8680 12238 8708 12406
rect 8864 12238 8892 12786
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10198 7052 10406
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6840 8430 6868 9862
rect 6932 9654 6960 10066
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6932 9178 6960 9590
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8090 6592 8230
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6472 7942 6592 7970
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6380 6730 6408 7822
rect 6472 7410 6500 7822
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5460 3602 5488 3946
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 4916 3292 5292 3301
rect 4972 3290 4996 3292
rect 5052 3290 5076 3292
rect 5132 3290 5156 3292
rect 5212 3290 5236 3292
rect 4972 3238 4982 3290
rect 5226 3238 5236 3290
rect 4972 3236 4996 3238
rect 5052 3236 5076 3238
rect 5132 3236 5156 3238
rect 5212 3236 5236 3238
rect 4916 3227 5292 3236
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4908 2650 4936 2994
rect 5552 2774 5580 3878
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5644 3194 5672 3674
rect 5828 3534 5856 4966
rect 6472 4162 6500 7210
rect 6564 6610 6592 7942
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6564 6582 6684 6610
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5234 6592 5578
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6656 5114 6684 6582
rect 6748 5234 6776 7346
rect 6840 5710 6868 8366
rect 6932 7954 6960 8774
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7024 7886 7052 8910
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7546 7052 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 7478 7144 10610
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 10062 7236 10542
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9586 7236 9998
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9110 7236 9522
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7300 8838 7328 10610
rect 7852 10130 7880 12106
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11898 8064 12038
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 8496 11150 8524 11698
rect 8588 11200 8616 12174
rect 9140 11762 9168 12786
rect 9232 12442 9260 13126
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11218 8984 11494
rect 9232 11370 9260 12378
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9140 11342 9260 11370
rect 8668 11212 8720 11218
rect 8588 11172 8668 11200
rect 8668 11154 8720 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 7932 11144 7984 11150
rect 8484 11144 8536 11150
rect 7932 11086 7984 11092
rect 8390 11112 8446 11121
rect 7944 10810 7972 11086
rect 8484 11086 8536 11092
rect 8390 11047 8446 11056
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 9722 7880 10066
rect 8404 9994 8432 11047
rect 8496 10674 8524 11086
rect 8680 10810 8708 11154
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10198 8616 10610
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8588 10062 8616 10134
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8498 7328 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 7954 7328 8434
rect 7392 8090 7420 9658
rect 8128 9654 8156 9930
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8220 9602 8248 9862
rect 8220 9574 8432 9602
rect 8404 9382 8432 9574
rect 8772 9382 8800 11018
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9518 8892 10406
rect 8956 10130 8984 11154
rect 9140 11150 9168 11342
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10810 9076 10950
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 8974 8248 9114
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8404 8906 8432 9318
rect 8496 8906 8524 9318
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8404 8498 8432 8842
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7208 6934 7236 7890
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 7206 7512 7822
rect 8404 7750 8432 8434
rect 8496 7886 8524 8842
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8090 8708 8774
rect 9048 8294 9076 10746
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 9217 9168 10474
rect 9232 10266 9260 11222
rect 9324 10588 9352 12106
rect 9416 11354 9444 13194
rect 9508 12986 9536 13330
rect 9692 12986 9720 13466
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9508 12850 9536 12922
rect 9784 12850 9812 13262
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9600 11898 9628 12106
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9876 11286 9904 13942
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 10674 9536 11154
rect 9772 11144 9824 11150
rect 9692 11104 9772 11132
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9404 10600 9456 10606
rect 9324 10560 9404 10588
rect 9404 10542 9456 10548
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9232 9602 9260 10202
rect 9416 9654 9444 10542
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9404 9648 9456 9654
rect 9232 9574 9352 9602
rect 9404 9590 9456 9596
rect 9126 9208 9182 9217
rect 9126 9143 9128 9152
rect 9180 9143 9182 9152
rect 9128 9114 9180 9120
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9048 7886 9076 8230
rect 9324 8090 9352 9574
rect 9508 9518 9536 9862
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 8974 9536 9454
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9600 8922 9628 9046
rect 9692 9042 9720 11104
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10810 9904 11086
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9968 10690 9996 13874
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12374 10088 12582
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 10152 12220 10180 13806
rect 10428 12434 10456 14214
rect 10520 14074 10548 14962
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10612 13705 10640 17064
rect 10916 15260 11292 15269
rect 10972 15258 10996 15260
rect 11052 15258 11076 15260
rect 11132 15258 11156 15260
rect 11212 15258 11236 15260
rect 10972 15206 10982 15258
rect 11226 15206 11236 15258
rect 10972 15204 10996 15206
rect 11052 15204 11076 15206
rect 11132 15204 11156 15206
rect 11212 15204 11236 15206
rect 10916 15195 11292 15204
rect 11716 15162 11744 17064
rect 12820 15162 12848 17064
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 13924 15026 13952 17064
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 13084 14816 13136 14822
rect 13728 14816 13780 14822
rect 13136 14776 13308 14804
rect 13084 14758 13136 14764
rect 10704 14346 10732 14758
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10916 14172 11292 14181
rect 10972 14170 10996 14172
rect 11052 14170 11076 14172
rect 11132 14170 11156 14172
rect 11212 14170 11236 14172
rect 10972 14118 10982 14170
rect 11226 14118 11236 14170
rect 10972 14116 10996 14118
rect 11052 14116 11076 14118
rect 11132 14116 11156 14118
rect 11212 14116 11236 14118
rect 10916 14107 11292 14116
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10598 13696 10654 13705
rect 10598 13631 10654 13640
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10336 12406 10456 12434
rect 10232 12232 10284 12238
rect 10152 12192 10232 12220
rect 10232 12174 10284 12180
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9784 10662 9996 10690
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9600 8894 9720 8922
rect 9586 8528 9642 8537
rect 9692 8514 9720 8894
rect 9784 8634 9812 10662
rect 10060 10554 10088 12038
rect 10244 11354 10272 12174
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10152 11150 10180 11222
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10140 10668 10192 10674
rect 10244 10656 10272 11290
rect 10192 10628 10272 10656
rect 10140 10610 10192 10616
rect 9968 10526 10088 10554
rect 9968 10470 9996 10526
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9382 9996 10406
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 8974 9996 9318
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9692 8486 9812 8514
rect 9586 8463 9588 8472
rect 9640 8463 9642 8472
rect 9588 8434 9640 8440
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7484 6798 7512 7142
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7760 6390 7788 7278
rect 7852 7206 7880 7686
rect 9324 7342 9352 8026
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 7002 7880 7142
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8404 7002 8432 7278
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6390 8064 6734
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 8404 6322 8432 6938
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 7852 5642 7880 6054
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6828 5160 6880 5166
rect 6656 5086 6776 5114
rect 6828 5102 6880 5108
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4468 6684 4966
rect 6748 4622 6776 5086
rect 6840 4622 6868 5102
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4480 6788 4486
rect 6656 4440 6736 4468
rect 6736 4422 6788 4428
rect 6748 4214 6776 4422
rect 6840 4282 6868 4558
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4282 7052 4422
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6736 4208 6788 4214
rect 6472 4146 6684 4162
rect 6736 4150 6788 4156
rect 6472 4140 6696 4146
rect 6472 4134 6644 4140
rect 6644 4082 6696 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3738 6408 3878
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5828 3126 5856 3470
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5920 3058 5948 3334
rect 6380 3194 6408 3402
rect 6932 3398 6960 4082
rect 7116 4078 7144 5510
rect 7852 5030 7880 5578
rect 8312 5302 8340 5646
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8404 5114 8432 5850
rect 8496 5846 8524 6394
rect 8588 6322 8616 7142
rect 9324 6798 9352 7278
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 9232 5914 9260 6666
rect 9416 5914 9444 7958
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9496 7472 9548 7478
rect 9600 7426 9628 7754
rect 9548 7420 9628 7426
rect 9496 7414 9628 7420
rect 9508 7398 9628 7414
rect 9692 7410 9720 7822
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6934 9536 7278
rect 9600 7002 9628 7398
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9784 7324 9812 8486
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9876 8090 9904 8434
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9968 7478 9996 8774
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10152 7750 10180 8502
rect 10336 8294 10364 12406
rect 10520 12356 10548 12718
rect 10704 12442 10732 14010
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11348 13326 11376 13874
rect 11440 13870 11468 14350
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 14074 11836 14214
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13530 11744 13738
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 10916 13084 11292 13093
rect 10972 13082 10996 13084
rect 11052 13082 11076 13084
rect 11132 13082 11156 13084
rect 11212 13082 11236 13084
rect 10972 13030 10982 13082
rect 11226 13030 11236 13082
rect 10972 13028 10996 13030
rect 11052 13028 11076 13030
rect 11132 13028 11156 13030
rect 11212 13028 11236 13030
rect 10916 13019 11292 13028
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10428 12328 10548 12356
rect 10428 12238 10456 12328
rect 10692 12300 10744 12306
rect 10612 12260 10692 12288
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11558 10456 12174
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10244 8266 10364 8294
rect 10244 8022 10272 8266
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9784 7296 9996 7324
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9600 6202 9628 6938
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9508 6174 9628 6202
rect 9784 6186 9812 6598
rect 9876 6390 9904 6938
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9772 6180 9824 6186
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 5370 9352 5646
rect 9508 5370 9536 6174
rect 9772 6122 9824 6128
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5846 9628 6054
rect 9784 5953 9812 6122
rect 9770 5944 9826 5953
rect 9770 5879 9826 5888
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 8404 5086 8524 5114
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8404 4214 8432 4966
rect 8496 4622 8524 5086
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7392 3738 7420 3878
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5552 2746 5672 2774
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5644 2446 5672 2746
rect 6012 2446 6040 3130
rect 6932 2446 6960 3334
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7116 2514 7144 3062
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7484 2446 7512 3334
rect 7852 3126 7880 3878
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 8404 3534 8432 4150
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 8588 2650 8616 4558
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8772 2446 8800 5306
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8864 4010 8892 4762
rect 9324 4758 9352 5306
rect 9600 5234 9628 5782
rect 9772 5704 9824 5710
rect 9770 5672 9772 5681
rect 9968 5692 9996 7296
rect 10152 7206 10180 7686
rect 10244 7478 10272 7958
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10060 6254 10088 7142
rect 10244 6798 10272 7414
rect 10336 7002 10364 8026
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6458 10272 6734
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10060 5778 10088 6190
rect 10244 6186 10272 6394
rect 10336 6254 10364 6938
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10244 5846 10272 6122
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9824 5672 9996 5692
rect 9826 5664 9996 5672
rect 9770 5607 9826 5616
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 4282 8984 4490
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9232 4146 9260 4558
rect 9324 4282 9352 4694
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9416 4214 9444 4422
rect 9784 4282 9812 5607
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9680 4208 9732 4214
rect 9864 4208 9916 4214
rect 9732 4156 9864 4162
rect 9680 4150 9916 4156
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9220 4140 9272 4146
rect 9692 4134 9904 4150
rect 9220 4082 9272 4088
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 9048 3534 9076 4082
rect 9128 4072 9180 4078
rect 9864 4072 9916 4078
rect 9678 4040 9734 4049
rect 9180 4020 9678 4026
rect 9128 4014 9678 4020
rect 9140 3998 9678 4014
rect 9916 4032 10088 4060
rect 10152 4049 10180 5714
rect 10428 5302 10456 11494
rect 10520 8820 10548 11562
rect 10612 8974 10640 12260
rect 10692 12242 10744 12248
rect 11244 12232 11296 12238
rect 11348 12220 11376 13262
rect 11440 12850 11468 13466
rect 11808 13326 11836 13874
rect 11992 13682 12020 14758
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 11900 13654 12020 13682
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11296 12192 11376 12220
rect 11244 12174 11296 12180
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11014 10732 12106
rect 10916 11996 11292 12005
rect 10972 11994 10996 11996
rect 11052 11994 11076 11996
rect 11132 11994 11156 11996
rect 11212 11994 11236 11996
rect 10972 11942 10982 11994
rect 11226 11942 11236 11994
rect 10972 11940 10996 11942
rect 11052 11940 11076 11942
rect 11132 11940 11156 11942
rect 11212 11940 11236 11942
rect 10916 11931 11292 11940
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11072 11150 11100 11698
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10810 10732 10950
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10796 9722 10824 11018
rect 11164 10996 11192 11698
rect 11348 11694 11376 12192
rect 11440 11898 11468 12786
rect 11808 12714 11836 13262
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10857 10968 11192 10996
rect 10857 10810 10885 10968
rect 10916 10908 11292 10917
rect 10972 10906 10996 10908
rect 11052 10906 11076 10908
rect 11132 10906 11156 10908
rect 11212 10906 11236 10908
rect 10972 10854 10982 10906
rect 11226 10854 11236 10906
rect 10972 10852 10996 10854
rect 11052 10852 11076 10854
rect 11132 10852 11156 10854
rect 11212 10852 11236 10854
rect 10916 10843 11292 10852
rect 10857 10804 10928 10810
rect 10857 10764 10876 10804
rect 10876 10746 10928 10752
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10266 10916 10406
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10876 10056 10928 10062
rect 10980 10044 11008 10678
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10928 10016 11008 10044
rect 10876 9998 10928 10004
rect 11072 9926 11100 10406
rect 11164 10198 11192 10746
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11348 10130 11376 11154
rect 11440 10674 11468 11834
rect 11532 10742 11560 12310
rect 11624 12306 11652 12582
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 10810 11652 11698
rect 11716 11218 11744 12174
rect 11808 12102 11836 12650
rect 11900 12434 11928 13654
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12986 12020 13262
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11980 12844 12032 12850
rect 12084 12832 12112 14214
rect 12176 14074 12204 14214
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12032 12804 12112 12832
rect 11980 12786 12032 12792
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11900 12406 12020 12434
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11830 11836 12038
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10736 11572 10742
rect 11572 10684 11652 10690
rect 11520 10678 11652 10684
rect 11428 10668 11480 10674
rect 11532 10662 11652 10678
rect 11808 10674 11836 11086
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11428 10610 11480 10616
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 10916 9820 11292 9829
rect 10972 9818 10996 9820
rect 11052 9818 11076 9820
rect 11132 9818 11156 9820
rect 11212 9818 11236 9820
rect 10972 9766 10982 9818
rect 11226 9766 11236 9818
rect 10972 9764 10996 9766
rect 11052 9764 11076 9766
rect 11132 9764 11156 9766
rect 11212 9764 11236 9766
rect 10916 9755 11292 9764
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 10704 8974 10732 9522
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10520 8792 10640 8820
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7546 10548 7686
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 5846 10640 8792
rect 10916 8732 11292 8741
rect 10972 8730 10996 8732
rect 11052 8730 11076 8732
rect 11132 8730 11156 8732
rect 11212 8730 11236 8732
rect 10972 8678 10982 8730
rect 11226 8678 11236 8730
rect 10972 8676 10996 8678
rect 11052 8676 11076 8678
rect 11132 8676 11156 8678
rect 11212 8676 11236 8678
rect 10916 8667 11292 8676
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 8022 11100 8366
rect 11348 8362 11376 9522
rect 11440 9110 11468 9862
rect 11532 9586 11560 9862
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 11624 8430 11652 10662
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11716 8566 11744 10610
rect 11900 9674 11928 10950
rect 11808 9646 11928 9674
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11612 8424 11664 8430
rect 11808 8412 11836 9646
rect 11900 9586 11928 9646
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11612 8366 11664 8372
rect 11716 8384 11836 8412
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7274 10732 7822
rect 10916 7644 11292 7653
rect 10972 7642 10996 7644
rect 11052 7642 11076 7644
rect 11132 7642 11156 7644
rect 11212 7642 11236 7644
rect 10972 7590 10982 7642
rect 11226 7590 11236 7642
rect 10972 7588 10996 7590
rect 11052 7588 11076 7590
rect 11132 7588 11156 7590
rect 11212 7588 11236 7590
rect 10916 7579 11292 7588
rect 11348 7478 11376 8298
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 6798 10732 7210
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 7002 11100 7142
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6322 10732 6734
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10796 5710 10824 6598
rect 10916 6556 11292 6565
rect 10972 6554 10996 6556
rect 11052 6554 11076 6556
rect 11132 6554 11156 6556
rect 11212 6554 11236 6556
rect 10972 6502 10982 6554
rect 11226 6502 11236 6554
rect 10972 6500 10996 6502
rect 11052 6500 11076 6502
rect 11132 6500 11156 6502
rect 11212 6500 11236 6502
rect 10916 6491 11292 6500
rect 11348 6458 11376 6666
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10980 5642 11008 6258
rect 11164 5914 11192 6258
rect 11716 6254 11744 8384
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11808 7206 11836 7822
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 6372 11836 7142
rect 11900 7002 11928 7822
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11808 6344 11928 6372
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5914 11652 6054
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11428 5704 11480 5710
rect 11716 5681 11744 6190
rect 11794 5944 11850 5953
rect 11794 5879 11796 5888
rect 11848 5879 11850 5888
rect 11796 5850 11848 5856
rect 11428 5646 11480 5652
rect 11702 5672 11758 5681
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10520 4554 10548 5578
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 9864 4014 9916 4020
rect 9678 3975 9734 3984
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3194 9076 3470
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9140 2774 9168 3878
rect 9784 3738 9812 3946
rect 10060 3942 10088 4032
rect 10138 4040 10194 4049
rect 10138 3975 10194 3984
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9140 2746 9352 2774
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9324 2378 9352 2746
rect 10336 2446 10364 4422
rect 10612 4078 10640 5578
rect 11440 5574 11468 5646
rect 11702 5607 11758 5616
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 10796 5234 10824 5510
rect 10916 5468 11292 5477
rect 10972 5466 10996 5468
rect 11052 5466 11076 5468
rect 11132 5466 11156 5468
rect 11212 5466 11236 5468
rect 10972 5414 10982 5466
rect 11226 5414 11236 5466
rect 10972 5412 10996 5414
rect 11052 5412 11076 5414
rect 11132 5412 11156 5414
rect 11212 5412 11236 5414
rect 10916 5403 11292 5412
rect 11808 5370 11836 5850
rect 11900 5642 11928 6344
rect 11992 5642 12020 12406
rect 12084 11898 12112 12582
rect 12176 12442 12204 13874
rect 12268 13530 12296 14350
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11626 12204 12378
rect 12256 11756 12308 11762
rect 12360 11744 12388 14214
rect 12636 14074 12664 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12728 13870 12756 14350
rect 12912 14278 12940 14758
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12452 12986 12480 13806
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12544 11762 12572 12310
rect 12308 11716 12388 11744
rect 12532 11756 12584 11762
rect 12256 11698 12308 11704
rect 12532 11698 12584 11704
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12268 10674 12296 11698
rect 12728 11014 12756 13806
rect 12912 13734 12940 14214
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 11694 12940 13670
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13096 12442 13124 12718
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13188 12374 13216 12718
rect 13280 12434 13308 14776
rect 13728 14758 13780 14764
rect 13740 14618 13768 14758
rect 13916 14716 14292 14725
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14156 14716
rect 14212 14714 14236 14716
rect 13972 14662 13982 14714
rect 14226 14662 14236 14714
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14156 14662
rect 14212 14660 14236 14662
rect 13916 14651 14292 14660
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13326 13860 13670
rect 13916 13628 14292 13637
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14156 13628
rect 14212 13626 14236 13628
rect 13972 13574 13982 13626
rect 14226 13574 14236 13626
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14156 13574
rect 14212 13572 14236 13574
rect 13916 13563 14292 13572
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12986 13860 13262
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13916 12540 14292 12549
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14156 12540
rect 14212 12538 14236 12540
rect 13972 12486 13982 12538
rect 14226 12486 14236 12538
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14156 12486
rect 14212 12484 14236 12486
rect 13916 12475 14292 12484
rect 13280 12406 13676 12434
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11898 13492 12106
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 13004 11354 13032 11766
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12544 10606 12572 10950
rect 13096 10742 13124 11494
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12176 9722 12204 9998
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 9722 12296 9862
rect 12360 9722 12388 9998
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12162 9208 12218 9217
rect 12162 9143 12218 9152
rect 12176 9110 12204 9143
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12360 8922 12388 9658
rect 12452 9586 12480 9930
rect 12820 9586 12848 10406
rect 13648 9994 13676 12406
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11762 13860 12242
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 10810 13860 11698
rect 13916 11452 14292 11461
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14156 11452
rect 14212 11450 14236 11452
rect 13972 11398 13982 11450
rect 14226 11398 14236 11450
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14156 11398
rect 14212 11396 14236 11398
rect 13916 11387 14292 11396
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10266 13768 10610
rect 13916 10364 14292 10373
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14156 10364
rect 14212 10362 14236 10364
rect 13972 10310 13982 10362
rect 14226 10310 14236 10362
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14156 10310
rect 14212 10308 14236 10310
rect 13916 10299 14292 10308
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 8974 12572 9454
rect 12820 9178 12848 9522
rect 13188 9382 13216 9930
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13372 9110 13400 9930
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 12268 8894 12388 8922
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12268 8634 12296 8894
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12360 8498 12388 8774
rect 12544 8498 12572 8910
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12636 8498 12664 8842
rect 13372 8566 13400 9046
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12624 8492 12676 8498
rect 12676 8452 12756 8480
rect 12624 8434 12676 8440
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12268 6662 12296 6938
rect 12636 6798 12664 7142
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12084 5914 12112 6190
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5681 12112 5714
rect 12070 5672 12126 5681
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11980 5636 12032 5642
rect 12070 5607 12126 5616
rect 11980 5578 12032 5584
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10980 5030 11008 5170
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10704 4146 10732 4966
rect 11900 4826 11928 5578
rect 12176 5234 12204 6598
rect 12636 6390 12664 6734
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12360 5710 12388 6190
rect 12636 5710 12664 6326
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12360 5234 12388 5646
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 10796 4554 10824 4762
rect 12268 4554 12296 4966
rect 12636 4622 12664 5646
rect 12728 5370 12756 8452
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5710 12848 6190
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12912 5370 12940 6122
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12728 5166 12756 5306
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 10916 4380 11292 4389
rect 10972 4378 10996 4380
rect 11052 4378 11076 4380
rect 11132 4378 11156 4380
rect 11212 4378 11236 4380
rect 10972 4326 10982 4378
rect 11226 4326 11236 4378
rect 10972 4324 10996 4326
rect 11052 4324 11076 4326
rect 11132 4324 11156 4326
rect 11212 4324 11236 4326
rect 10916 4315 11292 4324
rect 12452 4282 12480 4422
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10508 4072 10560 4078
rect 10414 4040 10470 4049
rect 10508 4014 10560 4020
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10414 3975 10470 3984
rect 10428 3194 10456 3975
rect 10520 3534 10548 4014
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10520 2650 10548 3470
rect 10612 3466 10640 3878
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10916 3292 11292 3301
rect 10972 3290 10996 3292
rect 11052 3290 11076 3292
rect 11132 3290 11156 3292
rect 11212 3290 11236 3292
rect 10972 3238 10982 3290
rect 11226 3238 11236 3290
rect 10972 3236 10996 3238
rect 11052 3236 11076 3238
rect 11132 3236 11156 3238
rect 11212 3236 11236 3238
rect 10916 3227 11292 3236
rect 12636 3058 12664 4558
rect 12808 4548 12860 4554
rect 12808 4490 12860 4496
rect 12820 4282 12848 4490
rect 13188 4282 13216 5170
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13556 4146 13584 5578
rect 13648 5370 13676 9930
rect 13916 9276 14292 9285
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14156 9276
rect 14212 9274 14236 9276
rect 13972 9222 13982 9274
rect 14226 9222 14236 9274
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14156 9222
rect 14212 9220 14236 9222
rect 13916 9211 14292 9220
rect 15028 8537 15056 17064
rect 15014 8528 15070 8537
rect 15014 8463 15070 8472
rect 13916 8188 14292 8197
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14156 8188
rect 14212 8186 14236 8188
rect 13972 8134 13982 8186
rect 14226 8134 14236 8186
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14156 8134
rect 14212 8132 14236 8134
rect 13916 8123 14292 8132
rect 13916 7100 14292 7109
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14156 7100
rect 14212 7098 14236 7100
rect 13972 7046 13982 7098
rect 14226 7046 14236 7098
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14156 7046
rect 14212 7044 14236 7046
rect 13916 7035 14292 7044
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13832 5574 13860 6394
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 13916 6012 14292 6021
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14156 6012
rect 14212 6010 14236 6012
rect 13972 5958 13982 6010
rect 14226 5958 14236 6010
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14156 5958
rect 14212 5956 14236 5958
rect 13916 5947 14292 5956
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13832 4486 13860 5170
rect 13916 4924 14292 4933
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14156 4924
rect 14212 4922 14236 4924
rect 13972 4870 13982 4922
rect 14226 4870 14236 4922
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14156 4870
rect 14212 4868 14236 4870
rect 13916 4859 14292 4868
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13916 3836 14292 3845
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14156 3836
rect 14212 3834 14236 3836
rect 13972 3782 13982 3834
rect 14226 3782 14236 3834
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14156 3782
rect 14212 3780 14236 3782
rect 13916 3771 14292 3780
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 11072 2514 11100 2790
rect 13464 2650 13492 2994
rect 13916 2748 14292 2757
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14156 2748
rect 14212 2746 14236 2748
rect 13972 2694 13982 2746
rect 14226 2694 14236 2746
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14156 2694
rect 14212 2692 14236 2694
rect 13916 2683 14292 2692
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 14384 2514 14412 4422
rect 14476 3194 14504 6190
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14568 2774 14596 5510
rect 14476 2746 14596 2774
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14476 2446 14504 2746
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 756 2304 808 2310
rect 756 2246 808 2252
rect 1952 2304 2004 2310
rect 3700 2304 3752 2310
rect 2004 2264 2084 2292
rect 1952 2246 2004 2252
rect 768 800 796 2246
rect 2056 800 2084 2264
rect 4712 2304 4764 2310
rect 3700 2246 3752 2252
rect 4632 2264 4712 2292
rect 3344 870 3464 898
rect 3344 800 3372 870
rect 754 0 810 800
rect 2042 0 2098 800
rect 3330 0 3386 800
rect 3436 762 3464 870
rect 3712 762 3740 2246
rect 4632 800 4660 2264
rect 6000 2304 6052 2310
rect 4712 2246 4764 2252
rect 5920 2264 6000 2292
rect 4916 2204 5292 2213
rect 4972 2202 4996 2204
rect 5052 2202 5076 2204
rect 5132 2202 5156 2204
rect 5212 2202 5236 2204
rect 4972 2150 4982 2202
rect 5226 2150 5236 2202
rect 4972 2148 4996 2150
rect 5052 2148 5076 2150
rect 5132 2148 5156 2150
rect 5212 2148 5236 2150
rect 4916 2139 5292 2148
rect 5920 800 5948 2264
rect 6000 2246 6052 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 7116 1170 7144 2246
rect 8680 1170 8708 2246
rect 7116 1142 7236 1170
rect 7208 800 7236 1142
rect 8496 1142 8708 1170
rect 8496 800 8524 1142
rect 9784 800 9812 2314
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 10916 2204 11292 2213
rect 10972 2202 10996 2204
rect 11052 2202 11076 2204
rect 11132 2202 11156 2204
rect 11212 2202 11236 2204
rect 10972 2150 10982 2202
rect 11226 2150 11236 2202
rect 10972 2148 10996 2150
rect 11052 2148 11076 2150
rect 11132 2148 11156 2150
rect 11212 2148 11236 2150
rect 10916 2139 11292 2148
rect 11072 870 11192 898
rect 11072 800 11100 870
rect 3436 734 3740 762
rect 4618 0 4674 800
rect 5906 0 5962 800
rect 7194 0 7250 800
rect 8482 0 8538 800
rect 9770 0 9826 800
rect 11058 0 11114 800
rect 11164 762 11192 870
rect 11348 762 11376 2246
rect 12360 800 12388 2246
rect 13740 1170 13768 2246
rect 13648 1142 13768 1170
rect 13648 800 13676 1142
rect 14936 800 14964 2314
rect 11164 734 11376 762
rect 12346 0 12402 800
rect 13634 0 13690 800
rect 14922 0 14978 800
<< via2 >>
rect 4916 15258 4972 15260
rect 4996 15258 5052 15260
rect 5076 15258 5132 15260
rect 5156 15258 5212 15260
rect 5236 15258 5292 15260
rect 4916 15206 4918 15258
rect 4918 15206 4970 15258
rect 4970 15206 4972 15258
rect 4996 15206 5034 15258
rect 5034 15206 5046 15258
rect 5046 15206 5052 15258
rect 5076 15206 5098 15258
rect 5098 15206 5110 15258
rect 5110 15206 5132 15258
rect 5156 15206 5162 15258
rect 5162 15206 5174 15258
rect 5174 15206 5212 15258
rect 5236 15206 5238 15258
rect 5238 15206 5290 15258
rect 5290 15206 5292 15258
rect 4916 15204 4972 15206
rect 4996 15204 5052 15206
rect 5076 15204 5132 15206
rect 5156 15204 5212 15206
rect 5236 15204 5292 15206
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 2226 13932 2282 13968
rect 2226 13912 2228 13932
rect 2228 13912 2280 13932
rect 2280 13912 2282 13932
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 3974 11600 4030 11656
rect 4916 14170 4972 14172
rect 4996 14170 5052 14172
rect 5076 14170 5132 14172
rect 5156 14170 5212 14172
rect 5236 14170 5292 14172
rect 4916 14118 4918 14170
rect 4918 14118 4970 14170
rect 4970 14118 4972 14170
rect 4996 14118 5034 14170
rect 5034 14118 5046 14170
rect 5046 14118 5052 14170
rect 5076 14118 5098 14170
rect 5098 14118 5110 14170
rect 5110 14118 5132 14170
rect 5156 14118 5162 14170
rect 5162 14118 5174 14170
rect 5174 14118 5212 14170
rect 5236 14118 5238 14170
rect 5238 14118 5290 14170
rect 5290 14118 5292 14170
rect 4916 14116 4972 14118
rect 4996 14116 5052 14118
rect 5076 14116 5132 14118
rect 5156 14116 5212 14118
rect 5236 14116 5292 14118
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 9218 13932 9274 13968
rect 9218 13912 9220 13932
rect 9220 13912 9272 13932
rect 9272 13912 9274 13932
rect 4916 13082 4972 13084
rect 4996 13082 5052 13084
rect 5076 13082 5132 13084
rect 5156 13082 5212 13084
rect 5236 13082 5292 13084
rect 4916 13030 4918 13082
rect 4918 13030 4970 13082
rect 4970 13030 4972 13082
rect 4996 13030 5034 13082
rect 5034 13030 5046 13082
rect 5046 13030 5052 13082
rect 5076 13030 5098 13082
rect 5098 13030 5110 13082
rect 5110 13030 5132 13082
rect 5156 13030 5162 13082
rect 5162 13030 5174 13082
rect 5174 13030 5212 13082
rect 5236 13030 5238 13082
rect 5238 13030 5290 13082
rect 5290 13030 5292 13082
rect 4916 13028 4972 13030
rect 4996 13028 5052 13030
rect 5076 13028 5132 13030
rect 5156 13028 5212 13030
rect 5236 13028 5292 13030
rect 4434 11756 4490 11792
rect 4434 11736 4436 11756
rect 4436 11736 4488 11756
rect 4488 11736 4490 11756
rect 4916 11994 4972 11996
rect 4996 11994 5052 11996
rect 5076 11994 5132 11996
rect 5156 11994 5212 11996
rect 5236 11994 5292 11996
rect 4916 11942 4918 11994
rect 4918 11942 4970 11994
rect 4970 11942 4972 11994
rect 4996 11942 5034 11994
rect 5034 11942 5046 11994
rect 5046 11942 5052 11994
rect 5076 11942 5098 11994
rect 5098 11942 5110 11994
rect 5110 11942 5132 11994
rect 5156 11942 5162 11994
rect 5162 11942 5174 11994
rect 5174 11942 5212 11994
rect 5236 11942 5238 11994
rect 5238 11942 5290 11994
rect 5290 11942 5292 11994
rect 4916 11940 4972 11942
rect 4996 11940 5052 11942
rect 5076 11940 5132 11942
rect 5156 11940 5212 11942
rect 5236 11940 5292 11942
rect 4894 11092 4896 11112
rect 4896 11092 4948 11112
rect 4948 11092 4950 11112
rect 4894 11056 4950 11092
rect 4916 10906 4972 10908
rect 4996 10906 5052 10908
rect 5076 10906 5132 10908
rect 5156 10906 5212 10908
rect 5236 10906 5292 10908
rect 4916 10854 4918 10906
rect 4918 10854 4970 10906
rect 4970 10854 4972 10906
rect 4996 10854 5034 10906
rect 5034 10854 5046 10906
rect 5046 10854 5052 10906
rect 5076 10854 5098 10906
rect 5098 10854 5110 10906
rect 5110 10854 5132 10906
rect 5156 10854 5162 10906
rect 5162 10854 5174 10906
rect 5174 10854 5212 10906
rect 5236 10854 5238 10906
rect 5238 10854 5290 10906
rect 5290 10854 5292 10906
rect 4916 10852 4972 10854
rect 4996 10852 5052 10854
rect 5076 10852 5132 10854
rect 5156 10852 5212 10854
rect 5236 10852 5292 10854
rect 4916 9818 4972 9820
rect 4996 9818 5052 9820
rect 5076 9818 5132 9820
rect 5156 9818 5212 9820
rect 5236 9818 5292 9820
rect 4916 9766 4918 9818
rect 4918 9766 4970 9818
rect 4970 9766 4972 9818
rect 4996 9766 5034 9818
rect 5034 9766 5046 9818
rect 5046 9766 5052 9818
rect 5076 9766 5098 9818
rect 5098 9766 5110 9818
rect 5110 9766 5132 9818
rect 5156 9766 5162 9818
rect 5162 9766 5174 9818
rect 5174 9766 5212 9818
rect 5236 9766 5238 9818
rect 5238 9766 5290 9818
rect 5290 9766 5292 9818
rect 4916 9764 4972 9766
rect 4996 9764 5052 9766
rect 5076 9764 5132 9766
rect 5156 9764 5212 9766
rect 5236 9764 5292 9766
rect 5722 11600 5778 11656
rect 5998 11736 6054 11792
rect 4916 8730 4972 8732
rect 4996 8730 5052 8732
rect 5076 8730 5132 8732
rect 5156 8730 5212 8732
rect 5236 8730 5292 8732
rect 4916 8678 4918 8730
rect 4918 8678 4970 8730
rect 4970 8678 4972 8730
rect 4996 8678 5034 8730
rect 5034 8678 5046 8730
rect 5046 8678 5052 8730
rect 5076 8678 5098 8730
rect 5098 8678 5110 8730
rect 5110 8678 5132 8730
rect 5156 8678 5162 8730
rect 5162 8678 5174 8730
rect 5174 8678 5212 8730
rect 5236 8678 5238 8730
rect 5238 8678 5290 8730
rect 5290 8678 5292 8730
rect 4916 8676 4972 8678
rect 4996 8676 5052 8678
rect 5076 8676 5132 8678
rect 5156 8676 5212 8678
rect 5236 8676 5292 8678
rect 4916 7642 4972 7644
rect 4996 7642 5052 7644
rect 5076 7642 5132 7644
rect 5156 7642 5212 7644
rect 5236 7642 5292 7644
rect 4916 7590 4918 7642
rect 4918 7590 4970 7642
rect 4970 7590 4972 7642
rect 4996 7590 5034 7642
rect 5034 7590 5046 7642
rect 5046 7590 5052 7642
rect 5076 7590 5098 7642
rect 5098 7590 5110 7642
rect 5110 7590 5132 7642
rect 5156 7590 5162 7642
rect 5162 7590 5174 7642
rect 5174 7590 5212 7642
rect 5236 7590 5238 7642
rect 5238 7590 5290 7642
rect 5290 7590 5292 7642
rect 4916 7588 4972 7590
rect 4996 7588 5052 7590
rect 5076 7588 5132 7590
rect 5156 7588 5212 7590
rect 5236 7588 5292 7590
rect 4916 6554 4972 6556
rect 4996 6554 5052 6556
rect 5076 6554 5132 6556
rect 5156 6554 5212 6556
rect 5236 6554 5292 6556
rect 4916 6502 4918 6554
rect 4918 6502 4970 6554
rect 4970 6502 4972 6554
rect 4996 6502 5034 6554
rect 5034 6502 5046 6554
rect 5046 6502 5052 6554
rect 5076 6502 5098 6554
rect 5098 6502 5110 6554
rect 5110 6502 5132 6554
rect 5156 6502 5162 6554
rect 5162 6502 5174 6554
rect 5174 6502 5212 6554
rect 5236 6502 5238 6554
rect 5238 6502 5290 6554
rect 5290 6502 5292 6554
rect 4916 6500 4972 6502
rect 4996 6500 5052 6502
rect 5076 6500 5132 6502
rect 5156 6500 5212 6502
rect 5236 6500 5292 6502
rect 4916 5466 4972 5468
rect 4996 5466 5052 5468
rect 5076 5466 5132 5468
rect 5156 5466 5212 5468
rect 5236 5466 5292 5468
rect 4916 5414 4918 5466
rect 4918 5414 4970 5466
rect 4970 5414 4972 5466
rect 4996 5414 5034 5466
rect 5034 5414 5046 5466
rect 5046 5414 5052 5466
rect 5076 5414 5098 5466
rect 5098 5414 5110 5466
rect 5110 5414 5132 5466
rect 5156 5414 5162 5466
rect 5162 5414 5174 5466
rect 5174 5414 5212 5466
rect 5236 5414 5238 5466
rect 5238 5414 5290 5466
rect 5290 5414 5292 5466
rect 4916 5412 4972 5414
rect 4996 5412 5052 5414
rect 5076 5412 5132 5414
rect 5156 5412 5212 5414
rect 5236 5412 5292 5414
rect 4916 4378 4972 4380
rect 4996 4378 5052 4380
rect 5076 4378 5132 4380
rect 5156 4378 5212 4380
rect 5236 4378 5292 4380
rect 4916 4326 4918 4378
rect 4918 4326 4970 4378
rect 4970 4326 4972 4378
rect 4996 4326 5034 4378
rect 5034 4326 5046 4378
rect 5046 4326 5052 4378
rect 5076 4326 5098 4378
rect 5098 4326 5110 4378
rect 5110 4326 5132 4378
rect 5156 4326 5162 4378
rect 5162 4326 5174 4378
rect 5174 4326 5212 4378
rect 5236 4326 5238 4378
rect 5238 4326 5290 4378
rect 5290 4326 5292 4378
rect 4916 4324 4972 4326
rect 4996 4324 5052 4326
rect 5076 4324 5132 4326
rect 5156 4324 5212 4326
rect 5236 4324 5292 4326
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 4916 3290 4972 3292
rect 4996 3290 5052 3292
rect 5076 3290 5132 3292
rect 5156 3290 5212 3292
rect 5236 3290 5292 3292
rect 4916 3238 4918 3290
rect 4918 3238 4970 3290
rect 4970 3238 4972 3290
rect 4996 3238 5034 3290
rect 5034 3238 5046 3290
rect 5046 3238 5052 3290
rect 5076 3238 5098 3290
rect 5098 3238 5110 3290
rect 5110 3238 5132 3290
rect 5156 3238 5162 3290
rect 5162 3238 5174 3290
rect 5174 3238 5212 3290
rect 5236 3238 5238 3290
rect 5238 3238 5290 3290
rect 5290 3238 5292 3290
rect 4916 3236 4972 3238
rect 4996 3236 5052 3238
rect 5076 3236 5132 3238
rect 5156 3236 5212 3238
rect 5236 3236 5292 3238
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 8390 11056 8446 11112
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 9126 9172 9182 9208
rect 9126 9152 9128 9172
rect 9128 9152 9180 9172
rect 9180 9152 9182 9172
rect 10916 15258 10972 15260
rect 10996 15258 11052 15260
rect 11076 15258 11132 15260
rect 11156 15258 11212 15260
rect 11236 15258 11292 15260
rect 10916 15206 10918 15258
rect 10918 15206 10970 15258
rect 10970 15206 10972 15258
rect 10996 15206 11034 15258
rect 11034 15206 11046 15258
rect 11046 15206 11052 15258
rect 11076 15206 11098 15258
rect 11098 15206 11110 15258
rect 11110 15206 11132 15258
rect 11156 15206 11162 15258
rect 11162 15206 11174 15258
rect 11174 15206 11212 15258
rect 11236 15206 11238 15258
rect 11238 15206 11290 15258
rect 11290 15206 11292 15258
rect 10916 15204 10972 15206
rect 10996 15204 11052 15206
rect 11076 15204 11132 15206
rect 11156 15204 11212 15206
rect 11236 15204 11292 15206
rect 10916 14170 10972 14172
rect 10996 14170 11052 14172
rect 11076 14170 11132 14172
rect 11156 14170 11212 14172
rect 11236 14170 11292 14172
rect 10916 14118 10918 14170
rect 10918 14118 10970 14170
rect 10970 14118 10972 14170
rect 10996 14118 11034 14170
rect 11034 14118 11046 14170
rect 11046 14118 11052 14170
rect 11076 14118 11098 14170
rect 11098 14118 11110 14170
rect 11110 14118 11132 14170
rect 11156 14118 11162 14170
rect 11162 14118 11174 14170
rect 11174 14118 11212 14170
rect 11236 14118 11238 14170
rect 11238 14118 11290 14170
rect 11290 14118 11292 14170
rect 10916 14116 10972 14118
rect 10996 14116 11052 14118
rect 11076 14116 11132 14118
rect 11156 14116 11212 14118
rect 11236 14116 11292 14118
rect 10598 13640 10654 13696
rect 9586 8492 9642 8528
rect 9586 8472 9588 8492
rect 9588 8472 9640 8492
rect 9640 8472 9642 8492
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 10916 13082 10972 13084
rect 10996 13082 11052 13084
rect 11076 13082 11132 13084
rect 11156 13082 11212 13084
rect 11236 13082 11292 13084
rect 10916 13030 10918 13082
rect 10918 13030 10970 13082
rect 10970 13030 10972 13082
rect 10996 13030 11034 13082
rect 11034 13030 11046 13082
rect 11046 13030 11052 13082
rect 11076 13030 11098 13082
rect 11098 13030 11110 13082
rect 11110 13030 11132 13082
rect 11156 13030 11162 13082
rect 11162 13030 11174 13082
rect 11174 13030 11212 13082
rect 11236 13030 11238 13082
rect 11238 13030 11290 13082
rect 11290 13030 11292 13082
rect 10916 13028 10972 13030
rect 10996 13028 11052 13030
rect 11076 13028 11132 13030
rect 11156 13028 11212 13030
rect 11236 13028 11292 13030
rect 9770 5888 9826 5944
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 9770 5652 9772 5672
rect 9772 5652 9824 5672
rect 9824 5652 9826 5672
rect 9770 5616 9826 5652
rect 9678 3984 9734 4040
rect 10916 11994 10972 11996
rect 10996 11994 11052 11996
rect 11076 11994 11132 11996
rect 11156 11994 11212 11996
rect 11236 11994 11292 11996
rect 10916 11942 10918 11994
rect 10918 11942 10970 11994
rect 10970 11942 10972 11994
rect 10996 11942 11034 11994
rect 11034 11942 11046 11994
rect 11046 11942 11052 11994
rect 11076 11942 11098 11994
rect 11098 11942 11110 11994
rect 11110 11942 11132 11994
rect 11156 11942 11162 11994
rect 11162 11942 11174 11994
rect 11174 11942 11212 11994
rect 11236 11942 11238 11994
rect 11238 11942 11290 11994
rect 11290 11942 11292 11994
rect 10916 11940 10972 11942
rect 10996 11940 11052 11942
rect 11076 11940 11132 11942
rect 11156 11940 11212 11942
rect 11236 11940 11292 11942
rect 10916 10906 10972 10908
rect 10996 10906 11052 10908
rect 11076 10906 11132 10908
rect 11156 10906 11212 10908
rect 11236 10906 11292 10908
rect 10916 10854 10918 10906
rect 10918 10854 10970 10906
rect 10970 10854 10972 10906
rect 10996 10854 11034 10906
rect 11034 10854 11046 10906
rect 11046 10854 11052 10906
rect 11076 10854 11098 10906
rect 11098 10854 11110 10906
rect 11110 10854 11132 10906
rect 11156 10854 11162 10906
rect 11162 10854 11174 10906
rect 11174 10854 11212 10906
rect 11236 10854 11238 10906
rect 11238 10854 11290 10906
rect 11290 10854 11292 10906
rect 10916 10852 10972 10854
rect 10996 10852 11052 10854
rect 11076 10852 11132 10854
rect 11156 10852 11212 10854
rect 11236 10852 11292 10854
rect 10916 9818 10972 9820
rect 10996 9818 11052 9820
rect 11076 9818 11132 9820
rect 11156 9818 11212 9820
rect 11236 9818 11292 9820
rect 10916 9766 10918 9818
rect 10918 9766 10970 9818
rect 10970 9766 10972 9818
rect 10996 9766 11034 9818
rect 11034 9766 11046 9818
rect 11046 9766 11052 9818
rect 11076 9766 11098 9818
rect 11098 9766 11110 9818
rect 11110 9766 11132 9818
rect 11156 9766 11162 9818
rect 11162 9766 11174 9818
rect 11174 9766 11212 9818
rect 11236 9766 11238 9818
rect 11238 9766 11290 9818
rect 11290 9766 11292 9818
rect 10916 9764 10972 9766
rect 10996 9764 11052 9766
rect 11076 9764 11132 9766
rect 11156 9764 11212 9766
rect 11236 9764 11292 9766
rect 10916 8730 10972 8732
rect 10996 8730 11052 8732
rect 11076 8730 11132 8732
rect 11156 8730 11212 8732
rect 11236 8730 11292 8732
rect 10916 8678 10918 8730
rect 10918 8678 10970 8730
rect 10970 8678 10972 8730
rect 10996 8678 11034 8730
rect 11034 8678 11046 8730
rect 11046 8678 11052 8730
rect 11076 8678 11098 8730
rect 11098 8678 11110 8730
rect 11110 8678 11132 8730
rect 11156 8678 11162 8730
rect 11162 8678 11174 8730
rect 11174 8678 11212 8730
rect 11236 8678 11238 8730
rect 11238 8678 11290 8730
rect 11290 8678 11292 8730
rect 10916 8676 10972 8678
rect 10996 8676 11052 8678
rect 11076 8676 11132 8678
rect 11156 8676 11212 8678
rect 11236 8676 11292 8678
rect 10916 7642 10972 7644
rect 10996 7642 11052 7644
rect 11076 7642 11132 7644
rect 11156 7642 11212 7644
rect 11236 7642 11292 7644
rect 10916 7590 10918 7642
rect 10918 7590 10970 7642
rect 10970 7590 10972 7642
rect 10996 7590 11034 7642
rect 11034 7590 11046 7642
rect 11046 7590 11052 7642
rect 11076 7590 11098 7642
rect 11098 7590 11110 7642
rect 11110 7590 11132 7642
rect 11156 7590 11162 7642
rect 11162 7590 11174 7642
rect 11174 7590 11212 7642
rect 11236 7590 11238 7642
rect 11238 7590 11290 7642
rect 11290 7590 11292 7642
rect 10916 7588 10972 7590
rect 10996 7588 11052 7590
rect 11076 7588 11132 7590
rect 11156 7588 11212 7590
rect 11236 7588 11292 7590
rect 10916 6554 10972 6556
rect 10996 6554 11052 6556
rect 11076 6554 11132 6556
rect 11156 6554 11212 6556
rect 11236 6554 11292 6556
rect 10916 6502 10918 6554
rect 10918 6502 10970 6554
rect 10970 6502 10972 6554
rect 10996 6502 11034 6554
rect 11034 6502 11046 6554
rect 11046 6502 11052 6554
rect 11076 6502 11098 6554
rect 11098 6502 11110 6554
rect 11110 6502 11132 6554
rect 11156 6502 11162 6554
rect 11162 6502 11174 6554
rect 11174 6502 11212 6554
rect 11236 6502 11238 6554
rect 11238 6502 11290 6554
rect 11290 6502 11292 6554
rect 10916 6500 10972 6502
rect 10996 6500 11052 6502
rect 11076 6500 11132 6502
rect 11156 6500 11212 6502
rect 11236 6500 11292 6502
rect 11794 5908 11850 5944
rect 11794 5888 11796 5908
rect 11796 5888 11848 5908
rect 11848 5888 11850 5908
rect 10138 3984 10194 4040
rect 11702 5616 11758 5672
rect 10916 5466 10972 5468
rect 10996 5466 11052 5468
rect 11076 5466 11132 5468
rect 11156 5466 11212 5468
rect 11236 5466 11292 5468
rect 10916 5414 10918 5466
rect 10918 5414 10970 5466
rect 10970 5414 10972 5466
rect 10996 5414 11034 5466
rect 11034 5414 11046 5466
rect 11046 5414 11052 5466
rect 11076 5414 11098 5466
rect 11098 5414 11110 5466
rect 11110 5414 11132 5466
rect 11156 5414 11162 5466
rect 11162 5414 11174 5466
rect 11174 5414 11212 5466
rect 11236 5414 11238 5466
rect 11238 5414 11290 5466
rect 11290 5414 11292 5466
rect 10916 5412 10972 5414
rect 10996 5412 11052 5414
rect 11076 5412 11132 5414
rect 11156 5412 11212 5414
rect 11236 5412 11292 5414
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 14156 14714 14212 14716
rect 14236 14714 14292 14716
rect 13916 14662 13918 14714
rect 13918 14662 13970 14714
rect 13970 14662 13972 14714
rect 13996 14662 14034 14714
rect 14034 14662 14046 14714
rect 14046 14662 14052 14714
rect 14076 14662 14098 14714
rect 14098 14662 14110 14714
rect 14110 14662 14132 14714
rect 14156 14662 14162 14714
rect 14162 14662 14174 14714
rect 14174 14662 14212 14714
rect 14236 14662 14238 14714
rect 14238 14662 14290 14714
rect 14290 14662 14292 14714
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 14156 14660 14212 14662
rect 14236 14660 14292 14662
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 14156 13626 14212 13628
rect 14236 13626 14292 13628
rect 13916 13574 13918 13626
rect 13918 13574 13970 13626
rect 13970 13574 13972 13626
rect 13996 13574 14034 13626
rect 14034 13574 14046 13626
rect 14046 13574 14052 13626
rect 14076 13574 14098 13626
rect 14098 13574 14110 13626
rect 14110 13574 14132 13626
rect 14156 13574 14162 13626
rect 14162 13574 14174 13626
rect 14174 13574 14212 13626
rect 14236 13574 14238 13626
rect 14238 13574 14290 13626
rect 14290 13574 14292 13626
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 14156 13572 14212 13574
rect 14236 13572 14292 13574
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 14156 12538 14212 12540
rect 14236 12538 14292 12540
rect 13916 12486 13918 12538
rect 13918 12486 13970 12538
rect 13970 12486 13972 12538
rect 13996 12486 14034 12538
rect 14034 12486 14046 12538
rect 14046 12486 14052 12538
rect 14076 12486 14098 12538
rect 14098 12486 14110 12538
rect 14110 12486 14132 12538
rect 14156 12486 14162 12538
rect 14162 12486 14174 12538
rect 14174 12486 14212 12538
rect 14236 12486 14238 12538
rect 14238 12486 14290 12538
rect 14290 12486 14292 12538
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 14156 12484 14212 12486
rect 14236 12484 14292 12486
rect 12162 9152 12218 9208
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 14156 11450 14212 11452
rect 14236 11450 14292 11452
rect 13916 11398 13918 11450
rect 13918 11398 13970 11450
rect 13970 11398 13972 11450
rect 13996 11398 14034 11450
rect 14034 11398 14046 11450
rect 14046 11398 14052 11450
rect 14076 11398 14098 11450
rect 14098 11398 14110 11450
rect 14110 11398 14132 11450
rect 14156 11398 14162 11450
rect 14162 11398 14174 11450
rect 14174 11398 14212 11450
rect 14236 11398 14238 11450
rect 14238 11398 14290 11450
rect 14290 11398 14292 11450
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 14156 11396 14212 11398
rect 14236 11396 14292 11398
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 14156 10362 14212 10364
rect 14236 10362 14292 10364
rect 13916 10310 13918 10362
rect 13918 10310 13970 10362
rect 13970 10310 13972 10362
rect 13996 10310 14034 10362
rect 14034 10310 14046 10362
rect 14046 10310 14052 10362
rect 14076 10310 14098 10362
rect 14098 10310 14110 10362
rect 14110 10310 14132 10362
rect 14156 10310 14162 10362
rect 14162 10310 14174 10362
rect 14174 10310 14212 10362
rect 14236 10310 14238 10362
rect 14238 10310 14290 10362
rect 14290 10310 14292 10362
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14156 10308 14212 10310
rect 14236 10308 14292 10310
rect 12070 5616 12126 5672
rect 10916 4378 10972 4380
rect 10996 4378 11052 4380
rect 11076 4378 11132 4380
rect 11156 4378 11212 4380
rect 11236 4378 11292 4380
rect 10916 4326 10918 4378
rect 10918 4326 10970 4378
rect 10970 4326 10972 4378
rect 10996 4326 11034 4378
rect 11034 4326 11046 4378
rect 11046 4326 11052 4378
rect 11076 4326 11098 4378
rect 11098 4326 11110 4378
rect 11110 4326 11132 4378
rect 11156 4326 11162 4378
rect 11162 4326 11174 4378
rect 11174 4326 11212 4378
rect 11236 4326 11238 4378
rect 11238 4326 11290 4378
rect 11290 4326 11292 4378
rect 10916 4324 10972 4326
rect 10996 4324 11052 4326
rect 11076 4324 11132 4326
rect 11156 4324 11212 4326
rect 11236 4324 11292 4326
rect 10414 3984 10470 4040
rect 10916 3290 10972 3292
rect 10996 3290 11052 3292
rect 11076 3290 11132 3292
rect 11156 3290 11212 3292
rect 11236 3290 11292 3292
rect 10916 3238 10918 3290
rect 10918 3238 10970 3290
rect 10970 3238 10972 3290
rect 10996 3238 11034 3290
rect 11034 3238 11046 3290
rect 11046 3238 11052 3290
rect 11076 3238 11098 3290
rect 11098 3238 11110 3290
rect 11110 3238 11132 3290
rect 11156 3238 11162 3290
rect 11162 3238 11174 3290
rect 11174 3238 11212 3290
rect 11236 3238 11238 3290
rect 11238 3238 11290 3290
rect 11290 3238 11292 3290
rect 10916 3236 10972 3238
rect 10996 3236 11052 3238
rect 11076 3236 11132 3238
rect 11156 3236 11212 3238
rect 11236 3236 11292 3238
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 14156 9274 14212 9276
rect 14236 9274 14292 9276
rect 13916 9222 13918 9274
rect 13918 9222 13970 9274
rect 13970 9222 13972 9274
rect 13996 9222 14034 9274
rect 14034 9222 14046 9274
rect 14046 9222 14052 9274
rect 14076 9222 14098 9274
rect 14098 9222 14110 9274
rect 14110 9222 14132 9274
rect 14156 9222 14162 9274
rect 14162 9222 14174 9274
rect 14174 9222 14212 9274
rect 14236 9222 14238 9274
rect 14238 9222 14290 9274
rect 14290 9222 14292 9274
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 14156 9220 14212 9222
rect 14236 9220 14292 9222
rect 15014 8472 15070 8528
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 14156 8186 14212 8188
rect 14236 8186 14292 8188
rect 13916 8134 13918 8186
rect 13918 8134 13970 8186
rect 13970 8134 13972 8186
rect 13996 8134 14034 8186
rect 14034 8134 14046 8186
rect 14046 8134 14052 8186
rect 14076 8134 14098 8186
rect 14098 8134 14110 8186
rect 14110 8134 14132 8186
rect 14156 8134 14162 8186
rect 14162 8134 14174 8186
rect 14174 8134 14212 8186
rect 14236 8134 14238 8186
rect 14238 8134 14290 8186
rect 14290 8134 14292 8186
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 14156 8132 14212 8134
rect 14236 8132 14292 8134
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 14156 7098 14212 7100
rect 14236 7098 14292 7100
rect 13916 7046 13918 7098
rect 13918 7046 13970 7098
rect 13970 7046 13972 7098
rect 13996 7046 14034 7098
rect 14034 7046 14046 7098
rect 14046 7046 14052 7098
rect 14076 7046 14098 7098
rect 14098 7046 14110 7098
rect 14110 7046 14132 7098
rect 14156 7046 14162 7098
rect 14162 7046 14174 7098
rect 14174 7046 14212 7098
rect 14236 7046 14238 7098
rect 14238 7046 14290 7098
rect 14290 7046 14292 7098
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14156 7044 14212 7046
rect 14236 7044 14292 7046
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 14156 6010 14212 6012
rect 14236 6010 14292 6012
rect 13916 5958 13918 6010
rect 13918 5958 13970 6010
rect 13970 5958 13972 6010
rect 13996 5958 14034 6010
rect 14034 5958 14046 6010
rect 14046 5958 14052 6010
rect 14076 5958 14098 6010
rect 14098 5958 14110 6010
rect 14110 5958 14132 6010
rect 14156 5958 14162 6010
rect 14162 5958 14174 6010
rect 14174 5958 14212 6010
rect 14236 5958 14238 6010
rect 14238 5958 14290 6010
rect 14290 5958 14292 6010
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14156 5956 14212 5958
rect 14236 5956 14292 5958
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 14156 4922 14212 4924
rect 14236 4922 14292 4924
rect 13916 4870 13918 4922
rect 13918 4870 13970 4922
rect 13970 4870 13972 4922
rect 13996 4870 14034 4922
rect 14034 4870 14046 4922
rect 14046 4870 14052 4922
rect 14076 4870 14098 4922
rect 14098 4870 14110 4922
rect 14110 4870 14132 4922
rect 14156 4870 14162 4922
rect 14162 4870 14174 4922
rect 14174 4870 14212 4922
rect 14236 4870 14238 4922
rect 14238 4870 14290 4922
rect 14290 4870 14292 4922
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14156 4868 14212 4870
rect 14236 4868 14292 4870
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 14156 3834 14212 3836
rect 14236 3834 14292 3836
rect 13916 3782 13918 3834
rect 13918 3782 13970 3834
rect 13970 3782 13972 3834
rect 13996 3782 14034 3834
rect 14034 3782 14046 3834
rect 14046 3782 14052 3834
rect 14076 3782 14098 3834
rect 14098 3782 14110 3834
rect 14110 3782 14132 3834
rect 14156 3782 14162 3834
rect 14162 3782 14174 3834
rect 14174 3782 14212 3834
rect 14236 3782 14238 3834
rect 14238 3782 14290 3834
rect 14290 3782 14292 3834
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14156 3780 14212 3782
rect 14236 3780 14292 3782
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 14156 2746 14212 2748
rect 14236 2746 14292 2748
rect 13916 2694 13918 2746
rect 13918 2694 13970 2746
rect 13970 2694 13972 2746
rect 13996 2694 14034 2746
rect 14034 2694 14046 2746
rect 14046 2694 14052 2746
rect 14076 2694 14098 2746
rect 14098 2694 14110 2746
rect 14110 2694 14132 2746
rect 14156 2694 14162 2746
rect 14162 2694 14174 2746
rect 14174 2694 14212 2746
rect 14236 2694 14238 2746
rect 14238 2694 14290 2746
rect 14290 2694 14292 2746
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 14156 2692 14212 2694
rect 14236 2692 14292 2694
rect 4916 2202 4972 2204
rect 4996 2202 5052 2204
rect 5076 2202 5132 2204
rect 5156 2202 5212 2204
rect 5236 2202 5292 2204
rect 4916 2150 4918 2202
rect 4918 2150 4970 2202
rect 4970 2150 4972 2202
rect 4996 2150 5034 2202
rect 5034 2150 5046 2202
rect 5046 2150 5052 2202
rect 5076 2150 5098 2202
rect 5098 2150 5110 2202
rect 5110 2150 5132 2202
rect 5156 2150 5162 2202
rect 5162 2150 5174 2202
rect 5174 2150 5212 2202
rect 5236 2150 5238 2202
rect 5238 2150 5290 2202
rect 5290 2150 5292 2202
rect 4916 2148 4972 2150
rect 4996 2148 5052 2150
rect 5076 2148 5132 2150
rect 5156 2148 5212 2150
rect 5236 2148 5292 2150
rect 10916 2202 10972 2204
rect 10996 2202 11052 2204
rect 11076 2202 11132 2204
rect 11156 2202 11212 2204
rect 11236 2202 11292 2204
rect 10916 2150 10918 2202
rect 10918 2150 10970 2202
rect 10970 2150 10972 2202
rect 10996 2150 11034 2202
rect 11034 2150 11046 2202
rect 11046 2150 11052 2202
rect 11076 2150 11098 2202
rect 11098 2150 11110 2202
rect 11110 2150 11132 2202
rect 11156 2150 11162 2202
rect 11162 2150 11174 2202
rect 11174 2150 11212 2202
rect 11236 2150 11238 2202
rect 11238 2150 11290 2202
rect 11290 2150 11292 2202
rect 10916 2148 10972 2150
rect 10996 2148 11052 2150
rect 11076 2148 11132 2150
rect 11156 2148 11212 2150
rect 11236 2148 11292 2150
<< metal3 >>
rect 4906 15264 5302 15265
rect 4906 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5072 15264
rect 5136 15200 5152 15264
rect 5216 15200 5232 15264
rect 5296 15200 5302 15264
rect 4906 15199 5302 15200
rect 10906 15264 11302 15265
rect 10906 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11072 15264
rect 11136 15200 11152 15264
rect 11216 15200 11232 15264
rect 11296 15200 11302 15264
rect 10906 15199 11302 15200
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 13906 14720 14302 14721
rect 13906 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14302 14720
rect 13906 14655 14302 14656
rect 4906 14176 5302 14177
rect 4906 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5302 14176
rect 4906 14111 5302 14112
rect 10906 14176 11302 14177
rect 10906 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11302 14176
rect 10906 14111 11302 14112
rect 2221 13970 2287 13973
rect 9213 13970 9279 13973
rect 2221 13968 9279 13970
rect 2221 13912 2226 13968
rect 2282 13912 9218 13968
rect 9274 13912 9279 13968
rect 2221 13910 9279 13912
rect 2221 13907 2287 13910
rect 9213 13907 9279 13910
rect 10593 13700 10659 13701
rect 10542 13698 10548 13700
rect 10502 13638 10548 13698
rect 10612 13696 10659 13700
rect 10654 13640 10659 13696
rect 10542 13636 10548 13638
rect 10612 13636 10659 13640
rect 10593 13635 10659 13636
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 13906 13632 14302 13633
rect 13906 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14302 13632
rect 13906 13567 14302 13568
rect 4906 13088 5302 13089
rect 4906 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5302 13088
rect 4906 13023 5302 13024
rect 10906 13088 11302 13089
rect 10906 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11302 13088
rect 10906 13023 11302 13024
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 13906 12544 14302 12545
rect 13906 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14302 12544
rect 13906 12479 14302 12480
rect 4906 12000 5302 12001
rect 4906 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5302 12000
rect 4906 11935 5302 11936
rect 10906 12000 11302 12001
rect 10906 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11302 12000
rect 10906 11935 11302 11936
rect 4429 11794 4495 11797
rect 5993 11794 6059 11797
rect 4429 11792 6059 11794
rect 4429 11736 4434 11792
rect 4490 11736 5998 11792
rect 6054 11736 6059 11792
rect 4429 11734 6059 11736
rect 4429 11731 4495 11734
rect 5993 11731 6059 11734
rect 3969 11658 4035 11661
rect 5717 11658 5783 11661
rect 3969 11656 5783 11658
rect 3969 11600 3974 11656
rect 4030 11600 5722 11656
rect 5778 11600 5783 11656
rect 3969 11598 5783 11600
rect 3969 11595 4035 11598
rect 5717 11595 5783 11598
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 13906 11456 14302 11457
rect 13906 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14302 11456
rect 13906 11391 14302 11392
rect 4889 11114 4955 11117
rect 8385 11114 8451 11117
rect 4889 11112 8451 11114
rect 4889 11056 4894 11112
rect 4950 11056 8390 11112
rect 8446 11056 8451 11112
rect 4889 11054 8451 11056
rect 4889 11051 4955 11054
rect 8385 11051 8451 11054
rect 4906 10912 5302 10913
rect 4906 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5302 10912
rect 4906 10847 5302 10848
rect 10906 10912 11302 10913
rect 10906 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11302 10912
rect 10906 10847 11302 10848
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 13906 10368 14302 10369
rect 13906 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14302 10368
rect 13906 10303 14302 10304
rect 4906 9824 5302 9825
rect 4906 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5302 9824
rect 4906 9759 5302 9760
rect 10906 9824 11302 9825
rect 10906 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11302 9824
rect 10906 9759 11302 9760
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 13906 9280 14302 9281
rect 13906 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14152 9280
rect 14216 9216 14232 9280
rect 14296 9216 14302 9280
rect 13906 9215 14302 9216
rect 9121 9210 9187 9213
rect 12157 9210 12223 9213
rect 9121 9208 12223 9210
rect 9121 9152 9126 9208
rect 9182 9152 12162 9208
rect 12218 9152 12223 9208
rect 9121 9150 12223 9152
rect 9121 9147 9187 9150
rect 12157 9147 12223 9150
rect 4906 8736 5302 8737
rect 4906 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5302 8736
rect 4906 8671 5302 8672
rect 10906 8736 11302 8737
rect 10906 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11302 8736
rect 10906 8671 11302 8672
rect 9581 8530 9647 8533
rect 15009 8530 15075 8533
rect 9581 8528 15075 8530
rect 9581 8472 9586 8528
rect 9642 8472 15014 8528
rect 15070 8472 15075 8528
rect 9581 8470 15075 8472
rect 9581 8467 9647 8470
rect 15009 8467 15075 8470
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 13906 8192 14302 8193
rect 13906 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14302 8192
rect 13906 8127 14302 8128
rect 4906 7648 5302 7649
rect 4906 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5302 7648
rect 4906 7583 5302 7584
rect 10906 7648 11302 7649
rect 10906 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11302 7648
rect 10906 7583 11302 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 13906 7104 14302 7105
rect 13906 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14302 7104
rect 13906 7039 14302 7040
rect 4906 6560 5302 6561
rect 4906 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5302 6560
rect 4906 6495 5302 6496
rect 10906 6560 11302 6561
rect 10906 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11302 6560
rect 10906 6495 11302 6496
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 13906 6016 14302 6017
rect 13906 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14302 6016
rect 13906 5951 14302 5952
rect 9765 5946 9831 5949
rect 11789 5946 11855 5949
rect 9765 5944 11855 5946
rect 9765 5888 9770 5944
rect 9826 5888 11794 5944
rect 11850 5888 11855 5944
rect 9765 5886 11855 5888
rect 9765 5883 9831 5886
rect 11789 5883 11855 5886
rect 9765 5674 9831 5677
rect 11697 5674 11763 5677
rect 12065 5674 12131 5677
rect 9765 5672 12131 5674
rect 9765 5616 9770 5672
rect 9826 5616 11702 5672
rect 11758 5616 12070 5672
rect 12126 5616 12131 5672
rect 9765 5614 12131 5616
rect 9765 5611 9831 5614
rect 11697 5611 11763 5614
rect 12065 5611 12131 5614
rect 4906 5472 5302 5473
rect 4906 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5302 5472
rect 4906 5407 5302 5408
rect 10906 5472 11302 5473
rect 10906 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11302 5472
rect 10906 5407 11302 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 13906 4928 14302 4929
rect 13906 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14302 4928
rect 13906 4863 14302 4864
rect 4906 4384 5302 4385
rect 4906 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5302 4384
rect 4906 4319 5302 4320
rect 10906 4384 11302 4385
rect 10906 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11302 4384
rect 10906 4319 11302 4320
rect 9673 4042 9739 4045
rect 10133 4042 10199 4045
rect 9673 4040 10199 4042
rect 9673 3984 9678 4040
rect 9734 3984 10138 4040
rect 10194 3984 10199 4040
rect 9673 3982 10199 3984
rect 9673 3979 9739 3982
rect 10133 3979 10199 3982
rect 10409 4042 10475 4045
rect 10542 4042 10548 4044
rect 10409 4040 10548 4042
rect 10409 3984 10414 4040
rect 10470 3984 10548 4040
rect 10409 3982 10548 3984
rect 10409 3979 10475 3982
rect 10542 3980 10548 3982
rect 10612 3980 10618 4044
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 13906 3840 14302 3841
rect 13906 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14302 3840
rect 13906 3775 14302 3776
rect 4906 3296 5302 3297
rect 4906 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5302 3296
rect 4906 3231 5302 3232
rect 10906 3296 11302 3297
rect 10906 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11302 3296
rect 10906 3231 11302 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 13906 2752 14302 2753
rect 13906 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14302 2752
rect 13906 2687 14302 2688
rect 4906 2208 5302 2209
rect 4906 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5302 2208
rect 4906 2143 5302 2144
rect 10906 2208 11302 2209
rect 10906 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11302 2208
rect 10906 2143 11302 2144
<< via3 >>
rect 4912 15260 4976 15264
rect 4912 15204 4916 15260
rect 4916 15204 4972 15260
rect 4972 15204 4976 15260
rect 4912 15200 4976 15204
rect 4992 15260 5056 15264
rect 4992 15204 4996 15260
rect 4996 15204 5052 15260
rect 5052 15204 5056 15260
rect 4992 15200 5056 15204
rect 5072 15260 5136 15264
rect 5072 15204 5076 15260
rect 5076 15204 5132 15260
rect 5132 15204 5136 15260
rect 5072 15200 5136 15204
rect 5152 15260 5216 15264
rect 5152 15204 5156 15260
rect 5156 15204 5212 15260
rect 5212 15204 5216 15260
rect 5152 15200 5216 15204
rect 5232 15260 5296 15264
rect 5232 15204 5236 15260
rect 5236 15204 5292 15260
rect 5292 15204 5296 15260
rect 5232 15200 5296 15204
rect 10912 15260 10976 15264
rect 10912 15204 10916 15260
rect 10916 15204 10972 15260
rect 10972 15204 10976 15260
rect 10912 15200 10976 15204
rect 10992 15260 11056 15264
rect 10992 15204 10996 15260
rect 10996 15204 11052 15260
rect 11052 15204 11056 15260
rect 10992 15200 11056 15204
rect 11072 15260 11136 15264
rect 11072 15204 11076 15260
rect 11076 15204 11132 15260
rect 11132 15204 11136 15260
rect 11072 15200 11136 15204
rect 11152 15260 11216 15264
rect 11152 15204 11156 15260
rect 11156 15204 11212 15260
rect 11212 15204 11216 15260
rect 11152 15200 11216 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 14152 14716 14216 14720
rect 14152 14660 14156 14716
rect 14156 14660 14212 14716
rect 14212 14660 14216 14716
rect 14152 14656 14216 14660
rect 14232 14716 14296 14720
rect 14232 14660 14236 14716
rect 14236 14660 14292 14716
rect 14292 14660 14296 14716
rect 14232 14656 14296 14660
rect 4912 14172 4976 14176
rect 4912 14116 4916 14172
rect 4916 14116 4972 14172
rect 4972 14116 4976 14172
rect 4912 14112 4976 14116
rect 4992 14172 5056 14176
rect 4992 14116 4996 14172
rect 4996 14116 5052 14172
rect 5052 14116 5056 14172
rect 4992 14112 5056 14116
rect 5072 14172 5136 14176
rect 5072 14116 5076 14172
rect 5076 14116 5132 14172
rect 5132 14116 5136 14172
rect 5072 14112 5136 14116
rect 5152 14172 5216 14176
rect 5152 14116 5156 14172
rect 5156 14116 5212 14172
rect 5212 14116 5216 14172
rect 5152 14112 5216 14116
rect 5232 14172 5296 14176
rect 5232 14116 5236 14172
rect 5236 14116 5292 14172
rect 5292 14116 5296 14172
rect 5232 14112 5296 14116
rect 10912 14172 10976 14176
rect 10912 14116 10916 14172
rect 10916 14116 10972 14172
rect 10972 14116 10976 14172
rect 10912 14112 10976 14116
rect 10992 14172 11056 14176
rect 10992 14116 10996 14172
rect 10996 14116 11052 14172
rect 11052 14116 11056 14172
rect 10992 14112 11056 14116
rect 11072 14172 11136 14176
rect 11072 14116 11076 14172
rect 11076 14116 11132 14172
rect 11132 14116 11136 14172
rect 11072 14112 11136 14116
rect 11152 14172 11216 14176
rect 11152 14116 11156 14172
rect 11156 14116 11212 14172
rect 11212 14116 11216 14172
rect 11152 14112 11216 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 10548 13696 10612 13700
rect 10548 13640 10598 13696
rect 10598 13640 10612 13696
rect 10548 13636 10612 13640
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 14152 13628 14216 13632
rect 14152 13572 14156 13628
rect 14156 13572 14212 13628
rect 14212 13572 14216 13628
rect 14152 13568 14216 13572
rect 14232 13628 14296 13632
rect 14232 13572 14236 13628
rect 14236 13572 14292 13628
rect 14292 13572 14296 13628
rect 14232 13568 14296 13572
rect 4912 13084 4976 13088
rect 4912 13028 4916 13084
rect 4916 13028 4972 13084
rect 4972 13028 4976 13084
rect 4912 13024 4976 13028
rect 4992 13084 5056 13088
rect 4992 13028 4996 13084
rect 4996 13028 5052 13084
rect 5052 13028 5056 13084
rect 4992 13024 5056 13028
rect 5072 13084 5136 13088
rect 5072 13028 5076 13084
rect 5076 13028 5132 13084
rect 5132 13028 5136 13084
rect 5072 13024 5136 13028
rect 5152 13084 5216 13088
rect 5152 13028 5156 13084
rect 5156 13028 5212 13084
rect 5212 13028 5216 13084
rect 5152 13024 5216 13028
rect 5232 13084 5296 13088
rect 5232 13028 5236 13084
rect 5236 13028 5292 13084
rect 5292 13028 5296 13084
rect 5232 13024 5296 13028
rect 10912 13084 10976 13088
rect 10912 13028 10916 13084
rect 10916 13028 10972 13084
rect 10972 13028 10976 13084
rect 10912 13024 10976 13028
rect 10992 13084 11056 13088
rect 10992 13028 10996 13084
rect 10996 13028 11052 13084
rect 11052 13028 11056 13084
rect 10992 13024 11056 13028
rect 11072 13084 11136 13088
rect 11072 13028 11076 13084
rect 11076 13028 11132 13084
rect 11132 13028 11136 13084
rect 11072 13024 11136 13028
rect 11152 13084 11216 13088
rect 11152 13028 11156 13084
rect 11156 13028 11212 13084
rect 11212 13028 11216 13084
rect 11152 13024 11216 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 14152 12540 14216 12544
rect 14152 12484 14156 12540
rect 14156 12484 14212 12540
rect 14212 12484 14216 12540
rect 14152 12480 14216 12484
rect 14232 12540 14296 12544
rect 14232 12484 14236 12540
rect 14236 12484 14292 12540
rect 14292 12484 14296 12540
rect 14232 12480 14296 12484
rect 4912 11996 4976 12000
rect 4912 11940 4916 11996
rect 4916 11940 4972 11996
rect 4972 11940 4976 11996
rect 4912 11936 4976 11940
rect 4992 11996 5056 12000
rect 4992 11940 4996 11996
rect 4996 11940 5052 11996
rect 5052 11940 5056 11996
rect 4992 11936 5056 11940
rect 5072 11996 5136 12000
rect 5072 11940 5076 11996
rect 5076 11940 5132 11996
rect 5132 11940 5136 11996
rect 5072 11936 5136 11940
rect 5152 11996 5216 12000
rect 5152 11940 5156 11996
rect 5156 11940 5212 11996
rect 5212 11940 5216 11996
rect 5152 11936 5216 11940
rect 5232 11996 5296 12000
rect 5232 11940 5236 11996
rect 5236 11940 5292 11996
rect 5292 11940 5296 11996
rect 5232 11936 5296 11940
rect 10912 11996 10976 12000
rect 10912 11940 10916 11996
rect 10916 11940 10972 11996
rect 10972 11940 10976 11996
rect 10912 11936 10976 11940
rect 10992 11996 11056 12000
rect 10992 11940 10996 11996
rect 10996 11940 11052 11996
rect 11052 11940 11056 11996
rect 10992 11936 11056 11940
rect 11072 11996 11136 12000
rect 11072 11940 11076 11996
rect 11076 11940 11132 11996
rect 11132 11940 11136 11996
rect 11072 11936 11136 11940
rect 11152 11996 11216 12000
rect 11152 11940 11156 11996
rect 11156 11940 11212 11996
rect 11212 11940 11216 11996
rect 11152 11936 11216 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 14152 11452 14216 11456
rect 14152 11396 14156 11452
rect 14156 11396 14212 11452
rect 14212 11396 14216 11452
rect 14152 11392 14216 11396
rect 14232 11452 14296 11456
rect 14232 11396 14236 11452
rect 14236 11396 14292 11452
rect 14292 11396 14296 11452
rect 14232 11392 14296 11396
rect 4912 10908 4976 10912
rect 4912 10852 4916 10908
rect 4916 10852 4972 10908
rect 4972 10852 4976 10908
rect 4912 10848 4976 10852
rect 4992 10908 5056 10912
rect 4992 10852 4996 10908
rect 4996 10852 5052 10908
rect 5052 10852 5056 10908
rect 4992 10848 5056 10852
rect 5072 10908 5136 10912
rect 5072 10852 5076 10908
rect 5076 10852 5132 10908
rect 5132 10852 5136 10908
rect 5072 10848 5136 10852
rect 5152 10908 5216 10912
rect 5152 10852 5156 10908
rect 5156 10852 5212 10908
rect 5212 10852 5216 10908
rect 5152 10848 5216 10852
rect 5232 10908 5296 10912
rect 5232 10852 5236 10908
rect 5236 10852 5292 10908
rect 5292 10852 5296 10908
rect 5232 10848 5296 10852
rect 10912 10908 10976 10912
rect 10912 10852 10916 10908
rect 10916 10852 10972 10908
rect 10972 10852 10976 10908
rect 10912 10848 10976 10852
rect 10992 10908 11056 10912
rect 10992 10852 10996 10908
rect 10996 10852 11052 10908
rect 11052 10852 11056 10908
rect 10992 10848 11056 10852
rect 11072 10908 11136 10912
rect 11072 10852 11076 10908
rect 11076 10852 11132 10908
rect 11132 10852 11136 10908
rect 11072 10848 11136 10852
rect 11152 10908 11216 10912
rect 11152 10852 11156 10908
rect 11156 10852 11212 10908
rect 11212 10852 11216 10908
rect 11152 10848 11216 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 14152 10364 14216 10368
rect 14152 10308 14156 10364
rect 14156 10308 14212 10364
rect 14212 10308 14216 10364
rect 14152 10304 14216 10308
rect 14232 10364 14296 10368
rect 14232 10308 14236 10364
rect 14236 10308 14292 10364
rect 14292 10308 14296 10364
rect 14232 10304 14296 10308
rect 4912 9820 4976 9824
rect 4912 9764 4916 9820
rect 4916 9764 4972 9820
rect 4972 9764 4976 9820
rect 4912 9760 4976 9764
rect 4992 9820 5056 9824
rect 4992 9764 4996 9820
rect 4996 9764 5052 9820
rect 5052 9764 5056 9820
rect 4992 9760 5056 9764
rect 5072 9820 5136 9824
rect 5072 9764 5076 9820
rect 5076 9764 5132 9820
rect 5132 9764 5136 9820
rect 5072 9760 5136 9764
rect 5152 9820 5216 9824
rect 5152 9764 5156 9820
rect 5156 9764 5212 9820
rect 5212 9764 5216 9820
rect 5152 9760 5216 9764
rect 5232 9820 5296 9824
rect 5232 9764 5236 9820
rect 5236 9764 5292 9820
rect 5292 9764 5296 9820
rect 5232 9760 5296 9764
rect 10912 9820 10976 9824
rect 10912 9764 10916 9820
rect 10916 9764 10972 9820
rect 10972 9764 10976 9820
rect 10912 9760 10976 9764
rect 10992 9820 11056 9824
rect 10992 9764 10996 9820
rect 10996 9764 11052 9820
rect 11052 9764 11056 9820
rect 10992 9760 11056 9764
rect 11072 9820 11136 9824
rect 11072 9764 11076 9820
rect 11076 9764 11132 9820
rect 11132 9764 11136 9820
rect 11072 9760 11136 9764
rect 11152 9820 11216 9824
rect 11152 9764 11156 9820
rect 11156 9764 11212 9820
rect 11212 9764 11216 9820
rect 11152 9760 11216 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 14152 9276 14216 9280
rect 14152 9220 14156 9276
rect 14156 9220 14212 9276
rect 14212 9220 14216 9276
rect 14152 9216 14216 9220
rect 14232 9276 14296 9280
rect 14232 9220 14236 9276
rect 14236 9220 14292 9276
rect 14292 9220 14296 9276
rect 14232 9216 14296 9220
rect 4912 8732 4976 8736
rect 4912 8676 4916 8732
rect 4916 8676 4972 8732
rect 4972 8676 4976 8732
rect 4912 8672 4976 8676
rect 4992 8732 5056 8736
rect 4992 8676 4996 8732
rect 4996 8676 5052 8732
rect 5052 8676 5056 8732
rect 4992 8672 5056 8676
rect 5072 8732 5136 8736
rect 5072 8676 5076 8732
rect 5076 8676 5132 8732
rect 5132 8676 5136 8732
rect 5072 8672 5136 8676
rect 5152 8732 5216 8736
rect 5152 8676 5156 8732
rect 5156 8676 5212 8732
rect 5212 8676 5216 8732
rect 5152 8672 5216 8676
rect 5232 8732 5296 8736
rect 5232 8676 5236 8732
rect 5236 8676 5292 8732
rect 5292 8676 5296 8732
rect 5232 8672 5296 8676
rect 10912 8732 10976 8736
rect 10912 8676 10916 8732
rect 10916 8676 10972 8732
rect 10972 8676 10976 8732
rect 10912 8672 10976 8676
rect 10992 8732 11056 8736
rect 10992 8676 10996 8732
rect 10996 8676 11052 8732
rect 11052 8676 11056 8732
rect 10992 8672 11056 8676
rect 11072 8732 11136 8736
rect 11072 8676 11076 8732
rect 11076 8676 11132 8732
rect 11132 8676 11136 8732
rect 11072 8672 11136 8676
rect 11152 8732 11216 8736
rect 11152 8676 11156 8732
rect 11156 8676 11212 8732
rect 11212 8676 11216 8732
rect 11152 8672 11216 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 14152 8188 14216 8192
rect 14152 8132 14156 8188
rect 14156 8132 14212 8188
rect 14212 8132 14216 8188
rect 14152 8128 14216 8132
rect 14232 8188 14296 8192
rect 14232 8132 14236 8188
rect 14236 8132 14292 8188
rect 14292 8132 14296 8188
rect 14232 8128 14296 8132
rect 4912 7644 4976 7648
rect 4912 7588 4916 7644
rect 4916 7588 4972 7644
rect 4972 7588 4976 7644
rect 4912 7584 4976 7588
rect 4992 7644 5056 7648
rect 4992 7588 4996 7644
rect 4996 7588 5052 7644
rect 5052 7588 5056 7644
rect 4992 7584 5056 7588
rect 5072 7644 5136 7648
rect 5072 7588 5076 7644
rect 5076 7588 5132 7644
rect 5132 7588 5136 7644
rect 5072 7584 5136 7588
rect 5152 7644 5216 7648
rect 5152 7588 5156 7644
rect 5156 7588 5212 7644
rect 5212 7588 5216 7644
rect 5152 7584 5216 7588
rect 5232 7644 5296 7648
rect 5232 7588 5236 7644
rect 5236 7588 5292 7644
rect 5292 7588 5296 7644
rect 5232 7584 5296 7588
rect 10912 7644 10976 7648
rect 10912 7588 10916 7644
rect 10916 7588 10972 7644
rect 10972 7588 10976 7644
rect 10912 7584 10976 7588
rect 10992 7644 11056 7648
rect 10992 7588 10996 7644
rect 10996 7588 11052 7644
rect 11052 7588 11056 7644
rect 10992 7584 11056 7588
rect 11072 7644 11136 7648
rect 11072 7588 11076 7644
rect 11076 7588 11132 7644
rect 11132 7588 11136 7644
rect 11072 7584 11136 7588
rect 11152 7644 11216 7648
rect 11152 7588 11156 7644
rect 11156 7588 11212 7644
rect 11212 7588 11216 7644
rect 11152 7584 11216 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 14152 7100 14216 7104
rect 14152 7044 14156 7100
rect 14156 7044 14212 7100
rect 14212 7044 14216 7100
rect 14152 7040 14216 7044
rect 14232 7100 14296 7104
rect 14232 7044 14236 7100
rect 14236 7044 14292 7100
rect 14292 7044 14296 7100
rect 14232 7040 14296 7044
rect 4912 6556 4976 6560
rect 4912 6500 4916 6556
rect 4916 6500 4972 6556
rect 4972 6500 4976 6556
rect 4912 6496 4976 6500
rect 4992 6556 5056 6560
rect 4992 6500 4996 6556
rect 4996 6500 5052 6556
rect 5052 6500 5056 6556
rect 4992 6496 5056 6500
rect 5072 6556 5136 6560
rect 5072 6500 5076 6556
rect 5076 6500 5132 6556
rect 5132 6500 5136 6556
rect 5072 6496 5136 6500
rect 5152 6556 5216 6560
rect 5152 6500 5156 6556
rect 5156 6500 5212 6556
rect 5212 6500 5216 6556
rect 5152 6496 5216 6500
rect 5232 6556 5296 6560
rect 5232 6500 5236 6556
rect 5236 6500 5292 6556
rect 5292 6500 5296 6556
rect 5232 6496 5296 6500
rect 10912 6556 10976 6560
rect 10912 6500 10916 6556
rect 10916 6500 10972 6556
rect 10972 6500 10976 6556
rect 10912 6496 10976 6500
rect 10992 6556 11056 6560
rect 10992 6500 10996 6556
rect 10996 6500 11052 6556
rect 11052 6500 11056 6556
rect 10992 6496 11056 6500
rect 11072 6556 11136 6560
rect 11072 6500 11076 6556
rect 11076 6500 11132 6556
rect 11132 6500 11136 6556
rect 11072 6496 11136 6500
rect 11152 6556 11216 6560
rect 11152 6500 11156 6556
rect 11156 6500 11212 6556
rect 11212 6500 11216 6556
rect 11152 6496 11216 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 14152 6012 14216 6016
rect 14152 5956 14156 6012
rect 14156 5956 14212 6012
rect 14212 5956 14216 6012
rect 14152 5952 14216 5956
rect 14232 6012 14296 6016
rect 14232 5956 14236 6012
rect 14236 5956 14292 6012
rect 14292 5956 14296 6012
rect 14232 5952 14296 5956
rect 4912 5468 4976 5472
rect 4912 5412 4916 5468
rect 4916 5412 4972 5468
rect 4972 5412 4976 5468
rect 4912 5408 4976 5412
rect 4992 5468 5056 5472
rect 4992 5412 4996 5468
rect 4996 5412 5052 5468
rect 5052 5412 5056 5468
rect 4992 5408 5056 5412
rect 5072 5468 5136 5472
rect 5072 5412 5076 5468
rect 5076 5412 5132 5468
rect 5132 5412 5136 5468
rect 5072 5408 5136 5412
rect 5152 5468 5216 5472
rect 5152 5412 5156 5468
rect 5156 5412 5212 5468
rect 5212 5412 5216 5468
rect 5152 5408 5216 5412
rect 5232 5468 5296 5472
rect 5232 5412 5236 5468
rect 5236 5412 5292 5468
rect 5292 5412 5296 5468
rect 5232 5408 5296 5412
rect 10912 5468 10976 5472
rect 10912 5412 10916 5468
rect 10916 5412 10972 5468
rect 10972 5412 10976 5468
rect 10912 5408 10976 5412
rect 10992 5468 11056 5472
rect 10992 5412 10996 5468
rect 10996 5412 11052 5468
rect 11052 5412 11056 5468
rect 10992 5408 11056 5412
rect 11072 5468 11136 5472
rect 11072 5412 11076 5468
rect 11076 5412 11132 5468
rect 11132 5412 11136 5468
rect 11072 5408 11136 5412
rect 11152 5468 11216 5472
rect 11152 5412 11156 5468
rect 11156 5412 11212 5468
rect 11212 5412 11216 5468
rect 11152 5408 11216 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 14152 4924 14216 4928
rect 14152 4868 14156 4924
rect 14156 4868 14212 4924
rect 14212 4868 14216 4924
rect 14152 4864 14216 4868
rect 14232 4924 14296 4928
rect 14232 4868 14236 4924
rect 14236 4868 14292 4924
rect 14292 4868 14296 4924
rect 14232 4864 14296 4868
rect 4912 4380 4976 4384
rect 4912 4324 4916 4380
rect 4916 4324 4972 4380
rect 4972 4324 4976 4380
rect 4912 4320 4976 4324
rect 4992 4380 5056 4384
rect 4992 4324 4996 4380
rect 4996 4324 5052 4380
rect 5052 4324 5056 4380
rect 4992 4320 5056 4324
rect 5072 4380 5136 4384
rect 5072 4324 5076 4380
rect 5076 4324 5132 4380
rect 5132 4324 5136 4380
rect 5072 4320 5136 4324
rect 5152 4380 5216 4384
rect 5152 4324 5156 4380
rect 5156 4324 5212 4380
rect 5212 4324 5216 4380
rect 5152 4320 5216 4324
rect 5232 4380 5296 4384
rect 5232 4324 5236 4380
rect 5236 4324 5292 4380
rect 5292 4324 5296 4380
rect 5232 4320 5296 4324
rect 10912 4380 10976 4384
rect 10912 4324 10916 4380
rect 10916 4324 10972 4380
rect 10972 4324 10976 4380
rect 10912 4320 10976 4324
rect 10992 4380 11056 4384
rect 10992 4324 10996 4380
rect 10996 4324 11052 4380
rect 11052 4324 11056 4380
rect 10992 4320 11056 4324
rect 11072 4380 11136 4384
rect 11072 4324 11076 4380
rect 11076 4324 11132 4380
rect 11132 4324 11136 4380
rect 11072 4320 11136 4324
rect 11152 4380 11216 4384
rect 11152 4324 11156 4380
rect 11156 4324 11212 4380
rect 11212 4324 11216 4380
rect 11152 4320 11216 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 10548 3980 10612 4044
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 14152 3836 14216 3840
rect 14152 3780 14156 3836
rect 14156 3780 14212 3836
rect 14212 3780 14216 3836
rect 14152 3776 14216 3780
rect 14232 3836 14296 3840
rect 14232 3780 14236 3836
rect 14236 3780 14292 3836
rect 14292 3780 14296 3836
rect 14232 3776 14296 3780
rect 4912 3292 4976 3296
rect 4912 3236 4916 3292
rect 4916 3236 4972 3292
rect 4972 3236 4976 3292
rect 4912 3232 4976 3236
rect 4992 3292 5056 3296
rect 4992 3236 4996 3292
rect 4996 3236 5052 3292
rect 5052 3236 5056 3292
rect 4992 3232 5056 3236
rect 5072 3292 5136 3296
rect 5072 3236 5076 3292
rect 5076 3236 5132 3292
rect 5132 3236 5136 3292
rect 5072 3232 5136 3236
rect 5152 3292 5216 3296
rect 5152 3236 5156 3292
rect 5156 3236 5212 3292
rect 5212 3236 5216 3292
rect 5152 3232 5216 3236
rect 5232 3292 5296 3296
rect 5232 3236 5236 3292
rect 5236 3236 5292 3292
rect 5292 3236 5296 3292
rect 5232 3232 5296 3236
rect 10912 3292 10976 3296
rect 10912 3236 10916 3292
rect 10916 3236 10972 3292
rect 10972 3236 10976 3292
rect 10912 3232 10976 3236
rect 10992 3292 11056 3296
rect 10992 3236 10996 3292
rect 10996 3236 11052 3292
rect 11052 3236 11056 3292
rect 10992 3232 11056 3236
rect 11072 3292 11136 3296
rect 11072 3236 11076 3292
rect 11076 3236 11132 3292
rect 11132 3236 11136 3292
rect 11072 3232 11136 3236
rect 11152 3292 11216 3296
rect 11152 3236 11156 3292
rect 11156 3236 11212 3292
rect 11212 3236 11216 3292
rect 11152 3232 11216 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 14152 2748 14216 2752
rect 14152 2692 14156 2748
rect 14156 2692 14212 2748
rect 14212 2692 14216 2748
rect 14152 2688 14216 2692
rect 14232 2748 14296 2752
rect 14232 2692 14236 2748
rect 14236 2692 14292 2748
rect 14292 2692 14296 2748
rect 14232 2688 14296 2692
rect 4912 2204 4976 2208
rect 4912 2148 4916 2204
rect 4916 2148 4972 2204
rect 4972 2148 4976 2204
rect 4912 2144 4976 2148
rect 4992 2204 5056 2208
rect 4992 2148 4996 2204
rect 4996 2148 5052 2204
rect 5052 2148 5056 2204
rect 4992 2144 5056 2148
rect 5072 2204 5136 2208
rect 5072 2148 5076 2204
rect 5076 2148 5132 2204
rect 5132 2148 5136 2204
rect 5072 2144 5136 2148
rect 5152 2204 5216 2208
rect 5152 2148 5156 2204
rect 5156 2148 5212 2204
rect 5212 2148 5216 2204
rect 5152 2144 5216 2148
rect 5232 2204 5296 2208
rect 5232 2148 5236 2204
rect 5236 2148 5292 2204
rect 5292 2148 5296 2204
rect 5232 2144 5296 2148
rect 10912 2204 10976 2208
rect 10912 2148 10916 2204
rect 10916 2148 10972 2204
rect 10972 2148 10976 2204
rect 10912 2144 10976 2148
rect 10992 2204 11056 2208
rect 10992 2148 10996 2204
rect 10996 2148 11052 2204
rect 11052 2148 11056 2204
rect 10992 2144 11056 2148
rect 11072 2204 11136 2208
rect 11072 2148 11076 2204
rect 11076 2148 11132 2204
rect 11132 2148 11136 2204
rect 11072 2144 11136 2148
rect 11152 2204 11216 2208
rect 11152 2148 11156 2204
rect 11156 2148 11212 2204
rect 11212 2148 11216 2204
rect 11152 2144 11216 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
<< metal4 >>
rect 1904 14720 2304 15280
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9280 2304 10304
rect 1904 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 8192 2304 9216
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 2752 2304 3776
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 4904 15264 5304 15280
rect 4904 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5072 15264
rect 5136 15200 5152 15264
rect 5216 15200 5232 15264
rect 5296 15200 5304 15264
rect 4904 14176 5304 15200
rect 4904 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5304 14176
rect 4904 13088 5304 14112
rect 4904 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5304 13088
rect 4904 12000 5304 13024
rect 4904 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5304 12000
rect 4904 10912 5304 11936
rect 4904 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5304 10912
rect 4904 9824 5304 10848
rect 4904 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5304 9824
rect 4904 8736 5304 9760
rect 4904 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5304 8736
rect 4904 7648 5304 8672
rect 4904 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5304 7648
rect 4904 6560 5304 7584
rect 4904 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5304 6560
rect 4904 5472 5304 6496
rect 4904 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5304 5472
rect 4904 4384 5304 5408
rect 4904 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5304 4384
rect 4904 3296 5304 4320
rect 4904 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5304 3296
rect 4904 2208 5304 3232
rect 4904 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5304 2208
rect 4904 2128 5304 2144
rect 7904 14720 8304 15280
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 10904 15264 11304 15280
rect 10904 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11072 15264
rect 11136 15200 11152 15264
rect 11216 15200 11232 15264
rect 11296 15200 11304 15264
rect 10904 14176 11304 15200
rect 10904 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11304 14176
rect 10547 13700 10613 13701
rect 10547 13636 10548 13700
rect 10612 13636 10613 13700
rect 10547 13635 10613 13636
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9280 8304 10304
rect 7904 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 8192 8304 9216
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 10550 4045 10610 13635
rect 10904 13088 11304 14112
rect 10904 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11304 13088
rect 10904 12000 11304 13024
rect 10904 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11304 12000
rect 10904 10912 11304 11936
rect 10904 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11304 10912
rect 10904 9824 11304 10848
rect 10904 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11304 9824
rect 10904 8736 11304 9760
rect 10904 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11304 8736
rect 10904 7648 11304 8672
rect 10904 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11304 7648
rect 10904 6560 11304 7584
rect 10904 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11304 6560
rect 10904 5472 11304 6496
rect 10904 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11304 5472
rect 10904 4384 11304 5408
rect 10904 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11304 4384
rect 10547 4044 10613 4045
rect 10547 3980 10548 4044
rect 10612 3980 10613 4044
rect 10547 3979 10613 3980
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 2752 8304 3776
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 10904 3296 11304 4320
rect 10904 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11304 3296
rect 10904 2208 11304 3232
rect 10904 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11304 2208
rect 10904 2128 11304 2144
rect 13904 14720 14304 15280
rect 13904 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14304 14720
rect 13904 13632 14304 14656
rect 13904 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14304 13632
rect 13904 12544 14304 13568
rect 13904 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14304 12544
rect 13904 11456 14304 12480
rect 13904 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14304 11456
rect 13904 10368 14304 11392
rect 13904 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14304 10368
rect 13904 9280 14304 10304
rect 13904 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14152 9280
rect 14216 9216 14232 9280
rect 14296 9216 14304 9280
rect 13904 8192 14304 9216
rect 13904 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14304 8192
rect 13904 7104 14304 8128
rect 13904 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14304 7104
rect 13904 6016 14304 7040
rect 13904 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14304 6016
rect 13904 4928 14304 5952
rect 13904 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14304 4928
rect 13904 3840 14304 4864
rect 13904 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14304 3840
rect 13904 2752 14304 3776
rect 13904 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14304 2752
rect 13904 2128 14304 2688
use sky130_fd_sc_hd__buf_2  _189_
timestamp 1713335925
transform -1 0 11500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_4  _190_
timestamp 1713335925
transform -1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _191_
timestamp 1713335925
transform -1 0 6256 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _192_
timestamp 1713335925
transform -1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp 1713335925
transform 1 0 11316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _194_
timestamp 1713335925
transform -1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1713335925
transform -1 0 8832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _196_
timestamp 1713335925
transform 1 0 10580 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _197_
timestamp 1713335925
transform -1 0 6164 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _198_
timestamp 1713335925
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _199_
timestamp 1713335925
transform -1 0 9660 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _200_
timestamp 1713335925
transform -1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _201_
timestamp 1713335925
transform -1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _202_
timestamp 1713335925
transform 1 0 5704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _203_
timestamp 1713335925
transform 1 0 7268 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _204_
timestamp 1713335925
transform 1 0 7820 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _205_
timestamp 1713335925
transform -1 0 9476 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _206_
timestamp 1713335925
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _207_
timestamp 1713335925
transform 1 0 7452 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _208_
timestamp 1713335925
transform -1 0 10856 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _209_
timestamp 1713335925
transform -1 0 8464 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _210_
timestamp 1713335925
transform -1 0 7912 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _211_
timestamp 1713335925
transform -1 0 4508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _212_
timestamp 1713335925
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1713335925
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _214_
timestamp 1713335925
transform 1 0 8648 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _215_
timestamp 1713335925
transform -1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1713335925
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _217_
timestamp 1713335925
transform -1 0 10672 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _218_
timestamp 1713335925
transform -1 0 13524 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _219_
timestamp 1713335925
transform 1 0 4600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1713335925
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _221_
timestamp 1713335925
transform 1 0 8556 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _222_
timestamp 1713335925
transform -1 0 8004 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _223_
timestamp 1713335925
transform 1 0 6992 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1713335925
transform 1 0 8280 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1713335925
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _226_
timestamp 1713335925
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1713335925
transform 1 0 6440 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _228_
timestamp 1713335925
transform -1 0 4692 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _229_
timestamp 1713335925
transform 1 0 6992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _230_
timestamp 1713335925
transform 1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _231_
timestamp 1713335925
transform 1 0 2576 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _232_
timestamp 1713335925
transform 1 0 2944 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _233_
timestamp 1713335925
transform 1 0 2024 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1713335925
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _235_
timestamp 1713335925
transform 1 0 5888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _236_
timestamp 1713335925
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _237_
timestamp 1713335925
transform 1 0 6532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _238_
timestamp 1713335925
transform -1 0 5888 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _239_
timestamp 1713335925
transform -1 0 5888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _240_
timestamp 1713335925
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _241_
timestamp 1713335925
transform 1 0 12788 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _242_
timestamp 1713335925
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _243_
timestamp 1713335925
transform -1 0 6992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _244_
timestamp 1713335925
transform 1 0 4600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1713335925
transform -1 0 7084 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _246_
timestamp 1713335925
transform 1 0 6440 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _247_
timestamp 1713335925
transform -1 0 6256 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _248_
timestamp 1713335925
transform 1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _249_
timestamp 1713335925
transform -1 0 10672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _250_
timestamp 1713335925
transform 1 0 12696 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _251_
timestamp 1713335925
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _252_
timestamp 1713335925
transform -1 0 13340 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _253_
timestamp 1713335925
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _254_
timestamp 1713335925
transform -1 0 6624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _255_
timestamp 1713335925
transform -1 0 6256 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _256_
timestamp 1713335925
transform -1 0 5060 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _257_
timestamp 1713335925
transform -1 0 8832 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _258_
timestamp 1713335925
transform -1 0 5888 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _259_
timestamp 1713335925
transform 1 0 4508 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _260_
timestamp 1713335925
transform 1 0 5060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _261_
timestamp 1713335925
transform -1 0 5428 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _262_
timestamp 1713335925
transform 1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _263_
timestamp 1713335925
transform 1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _264_
timestamp 1713335925
transform -1 0 5704 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _265_
timestamp 1713335925
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _266_
timestamp 1713335925
transform 1 0 2944 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp 1713335925
transform -1 0 5428 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _268_
timestamp 1713335925
transform -1 0 4968 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _269_
timestamp 1713335925
transform -1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _270_
timestamp 1713335925
transform -1 0 2760 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1713335925
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _272_
timestamp 1713335925
transform 1 0 3772 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _273_
timestamp 1713335925
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _274_
timestamp 1713335925
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _275_
timestamp 1713335925
transform 1 0 2944 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _276_
timestamp 1713335925
transform -1 0 2208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1713335925
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 1713335925
transform 1 0 12144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _279_
timestamp 1713335925
transform 1 0 9476 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1713335925
transform 1 0 9568 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _281_
timestamp 1713335925
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _282_
timestamp 1713335925
transform 1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1713335925
transform -1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _284_
timestamp 1713335925
transform 1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _285_
timestamp 1713335925
transform -1 0 12788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _286_
timestamp 1713335925
transform -1 0 8740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _287_
timestamp 1713335925
transform -1 0 8832 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _288_
timestamp 1713335925
transform 1 0 9016 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1713335925
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1713335925
transform -1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _291_
timestamp 1713335925
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _292_
timestamp 1713335925
transform 1 0 10948 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _293_
timestamp 1713335925
transform 1 0 13340 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _294_
timestamp 1713335925
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _295_
timestamp 1713335925
transform -1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _296_
timestamp 1713335925
transform 1 0 9384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _297_
timestamp 1713335925
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _298_
timestamp 1713335925
transform 1 0 10120 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _299_
timestamp 1713335925
transform 1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1713335925
transform 1 0 11040 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _301_
timestamp 1713335925
transform -1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _302_
timestamp 1713335925
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _303_
timestamp 1713335925
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _304_
timestamp 1713335925
transform -1 0 10580 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1713335925
transform -1 0 13984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _306_
timestamp 1713335925
transform 1 0 11500 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp 1713335925
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _308_
timestamp 1713335925
transform -1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _309_
timestamp 1713335925
transform -1 0 12512 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _310_
timestamp 1713335925
transform 1 0 12236 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _311_
timestamp 1713335925
transform -1 0 13616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _312_
timestamp 1713335925
transform 1 0 11776 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _313_
timestamp 1713335925
transform -1 0 12788 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1713335925
transform 1 0 13248 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _315_
timestamp 1713335925
transform -1 0 13616 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _316_
timestamp 1713335925
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _317_
timestamp 1713335925
transform -1 0 8096 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _318_
timestamp 1713335925
transform 1 0 8096 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _319_
timestamp 1713335925
transform -1 0 7728 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _320_
timestamp 1713335925
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _321_
timestamp 1713335925
transform -1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _322_
timestamp 1713335925
transform -1 0 3864 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1713335925
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _324_
timestamp 1713335925
transform 1 0 3220 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _325_
timestamp 1713335925
transform -1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1713335925
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _327_
timestamp 1713335925
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 1713335925
transform -1 0 3680 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1713335925
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _330_
timestamp 1713335925
transform 1 0 4232 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _331_
timestamp 1713335925
transform -1 0 4876 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1713335925
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _333_
timestamp 1713335925
transform 1 0 4876 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _334_
timestamp 1713335925
transform -1 0 5980 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1713335925
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _336_
timestamp 1713335925
transform -1 0 6992 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _337_
timestamp 1713335925
transform 1 0 5520 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1713335925
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _339_
timestamp 1713335925
transform 1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 1713335925
transform 1 0 5336 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1713335925
transform -1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _342_
timestamp 1713335925
transform 1 0 6440 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1713335925
transform 1 0 6992 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1713335925
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _345_
timestamp 1713335925
transform 1 0 7636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _346_
timestamp 1713335925
transform 1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _347_
timestamp 1713335925
transform 1 0 10672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _348_
timestamp 1713335925
transform -1 0 11040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _349_
timestamp 1713335925
transform 1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _350_
timestamp 1713335925
transform 1 0 10028 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _351_
timestamp 1713335925
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _352_
timestamp 1713335925
transform -1 0 11224 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _353_
timestamp 1713335925
transform -1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _354_
timestamp 1713335925
transform 1 0 9292 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _355_
timestamp 1713335925
transform 1 0 9844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _356_
timestamp 1713335925
transform 1 0 7820 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _357_
timestamp 1713335925
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _358_
timestamp 1713335925
transform -1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _359_
timestamp 1713335925
transform 1 0 11868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _360_
timestamp 1713335925
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _361_
timestamp 1713335925
transform -1 0 14076 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _362_
timestamp 1713335925
transform 1 0 11868 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _363_
timestamp 1713335925
transform 1 0 12052 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1713335925
transform -1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1713335925
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _366_
timestamp 1713335925
transform -1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _367_
timestamp 1713335925
transform -1 0 8464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _368_
timestamp 1713335925
transform -1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _369_
timestamp 1713335925
transform 1 0 9844 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _370_
timestamp 1713335925
transform 1 0 9108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _371_
timestamp 1713335925
transform 1 0 8556 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _372_
timestamp 1713335925
transform 1 0 4600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _373_
timestamp 1713335925
transform 1 0 3496 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _374_
timestamp 1713335925
transform 1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _375_
timestamp 1713335925
transform 1 0 2300 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _376_
timestamp 1713335925
transform -1 0 2300 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1713335925
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1713335925
transform 1 0 2024 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1713335925
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1713335925
transform 1 0 6624 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1713335925
transform 1 0 5152 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1713335925
transform 1 0 3588 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1713335925
transform -1 0 13984 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1713335925
transform 1 0 1840 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1713335925
transform 1 0 1380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1713335925
transform 1 0 12604 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1713335925
transform 1 0 12788 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1713335925
transform 1 0 9844 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1713335925
transform -1 0 8832 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1713335925
transform 1 0 10580 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _391_
timestamp 1713335925
transform 1 0 12512 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1713335925
transform 1 0 12696 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1713335925
transform 1 0 1932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1713335925
transform 1 0 1564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1713335925
transform 1 0 2208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1713335925
transform 1 0 3128 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1713335925
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1713335925
transform 1 0 5980 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1713335925
transform -1 0 6256 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1713335925
transform 1 0 7176 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1713335925
transform 1 0 11500 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _402_
timestamp 1713335925
transform 1 0 10396 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _403_
timestamp 1713335925
transform 1 0 5888 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _404_
timestamp 1713335925
transform 1 0 9016 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1713335925
transform 1 0 12512 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1713335925
transform 1 0 12512 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1713335925
transform 1 0 7728 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1713335925
transform 1 0 9200 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1713335925
transform -1 0 8832 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1713335925
transform 1 0 1380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1713335925
transform -1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1713335925
transform -1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1713335925
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1713335925
transform -1 0 6900 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1713335925
transform -1 0 6440 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1713335925
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1713335925
transform 1 0 10764 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_6
timestamp 1713335925
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_35
timestamp 1713335925
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45
timestamp 1713335925
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57
timestamp 1713335925
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1713335925
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_107
timestamp 1713335925
transform 1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1713335925
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_121
timestamp 1713335925
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_126
timestamp 1713335925
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1713335925
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1713335925
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_15
timestamp 1713335925
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 1713335925
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1713335925
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_60
timestamp 1713335925
transform 1 0 6624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_88
timestamp 1713335925
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_102
timestamp 1713335925
transform 1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107
timestamp 1713335925
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1713335925
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1713335925
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_141
timestamp 1713335925
transform 1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1713335925
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_15
timestamp 1713335925
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_20
timestamp 1713335925
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 1713335925
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 1713335925
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1713335925
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1713335925
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1713335925
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1713335925
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_95
timestamp 1713335925
transform 1 0 9844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_107
timestamp 1713335925
transform 1 0 10948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_119
timestamp 1713335925
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_131
timestamp 1713335925
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1713335925
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1713335925
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 1713335925
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_9
timestamp 1713335925
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_13
timestamp 1713335925
transform 1 0 2300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_21
timestamp 1713335925
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_28
timestamp 1713335925
transform 1 0 3680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1713335925
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_69
timestamp 1713335925
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_73
timestamp 1713335925
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_80
timestamp 1713335925
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_100
timestamp 1713335925
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_108
timestamp 1713335925
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1713335925
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_128
timestamp 1713335925
transform 1 0 12880 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_134
timestamp 1713335925
transform 1 0 13432 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_138
timestamp 1713335925
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_142
timestamp 1713335925
transform 1 0 14168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1713335925
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1713335925
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1713335925
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_36
timestamp 1713335925
transform 1 0 4416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_48
timestamp 1713335925
transform 1 0 5520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_56
timestamp 1713335925
transform 1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1713335925
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1713335925
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1713335925
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_89
timestamp 1713335925
transform 1 0 9292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_118
timestamp 1713335925
transform 1 0 11960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1713335925
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1713335925
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_15
timestamp 1713335925
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_35
timestamp 1713335925
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_39
timestamp 1713335925
transform 1 0 4692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_62
timestamp 1713335925
transform 1 0 6808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_70
timestamp 1713335925
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_78
timestamp 1713335925
transform 1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_84
timestamp 1713335925
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_88
timestamp 1713335925
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_100
timestamp 1713335925
transform 1 0 10304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1713335925
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1713335925
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1713335925
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_124
timestamp 1713335925
transform 1 0 12512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_141
timestamp 1713335925
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1713335925
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_11
timestamp 1713335925
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_17
timestamp 1713335925
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1713335925
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_72
timestamp 1713335925
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1713335925
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85
timestamp 1713335925
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_94
timestamp 1713335925
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_101
timestamp 1713335925
transform 1 0 10396 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_109
timestamp 1713335925
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_123
timestamp 1713335925
transform 1 0 12420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1713335925
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1713335925
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_30
timestamp 1713335925
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_38
timestamp 1713335925
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1713335925
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1713335925
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_69
timestamp 1713335925
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_84
timestamp 1713335925
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_92
timestamp 1713335925
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1713335925
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1713335925
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_140
timestamp 1713335925
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1713335925
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1713335925
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1713335925
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_69
timestamp 1713335925
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_75
timestamp 1713335925
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1713335925
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_104
timestamp 1713335925
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_108
timestamp 1713335925
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_129
timestamp 1713335925
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1713335925
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1713335925
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1713335925
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1713335925
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_23
timestamp 1713335925
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1713335925
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_42
timestamp 1713335925
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_48
timestamp 1713335925
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1713335925
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_90
timestamp 1713335925
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_96
timestamp 1713335925
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1713335925
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_133
timestamp 1713335925
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_141
timestamp 1713335925
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1713335925
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1713335925
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1713335925
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_36
timestamp 1713335925
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_63
timestamp 1713335925
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_73
timestamp 1713335925
transform 1 0 7820 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1713335925
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_91
timestamp 1713335925
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_122
timestamp 1713335925
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1713335925
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1713335925
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 1713335925
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_11
timestamp 1713335925
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_16
timestamp 1713335925
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_28
timestamp 1713335925
transform 1 0 3680 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_40
timestamp 1713335925
transform 1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1713335925
transform 1 0 5336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1713335925
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_60
timestamp 1713335925
transform 1 0 6624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_72
timestamp 1713335925
transform 1 0 7728 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_99
timestamp 1713335925
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1713335925
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_113
timestamp 1713335925
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_119
timestamp 1713335925
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_131
timestamp 1713335925
transform 1 0 13156 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1713335925
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1713335925
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1713335925
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1713335925
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_39
timestamp 1713335925
transform 1 0 4692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_47
timestamp 1713335925
transform 1 0 5428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_55
timestamp 1713335925
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_70
timestamp 1713335925
transform 1 0 7544 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1713335925
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_115
timestamp 1713335925
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_119
timestamp 1713335925
transform 1 0 12052 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1713335925
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1713335925
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1713335925
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1713335925
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_10
timestamp 1713335925
transform 1 0 2024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_18
timestamp 1713335925
transform 1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_27
timestamp 1713335925
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1713335925
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1713335925
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_64
timestamp 1713335925
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_70
timestamp 1713335925
transform 1 0 7544 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_91
timestamp 1713335925
transform 1 0 9476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_99
timestamp 1713335925
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1713335925
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_117
timestamp 1713335925
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1713335925
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1713335925
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_74
timestamp 1713335925
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_80
timestamp 1713335925
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1713335925
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_97
timestamp 1713335925
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_105
timestamp 1713335925
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_110
timestamp 1713335925
transform 1 0 11224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_118
timestamp 1713335925
transform 1 0 11960 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_123
timestamp 1713335925
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1713335925
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1713335925
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1713335925
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_19
timestamp 1713335925
transform 1 0 2852 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_25
timestamp 1713335925
transform 1 0 3404 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_35
timestamp 1713335925
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_50
timestamp 1713335925
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1713335925
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_65
timestamp 1713335925
transform 1 0 7084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_77
timestamp 1713335925
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_81
timestamp 1713335925
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_88
timestamp 1713335925
transform 1 0 9200 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_104
timestamp 1713335925
transform 1 0 10672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_120
timestamp 1713335925
transform 1 0 12144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_141
timestamp 1713335925
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1713335925
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_20
timestamp 1713335925
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_46
timestamp 1713335925
transform 1 0 5336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_65
timestamp 1713335925
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 1713335925
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_98
timestamp 1713335925
transform 1 0 10120 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_104
timestamp 1713335925
transform 1 0 10672 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_125
timestamp 1713335925
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1713335925
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1713335925
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1713335925
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1713335925
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_27
timestamp 1713335925
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_34
timestamp 1713335925
transform 1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1713335925
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1713335925
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1713335925
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_85
timestamp 1713335925
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_97
timestamp 1713335925
transform 1 0 10028 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_103
timestamp 1713335925
transform 1 0 10580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_118
timestamp 1713335925
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_136
timestamp 1713335925
transform 1 0 13616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_142
timestamp 1713335925
transform 1 0 14168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 1713335925
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1713335925
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 1713335925
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1713335925
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_43
timestamp 1713335925
transform 1 0 5060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_56
timestamp 1713335925
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_65
timestamp 1713335925
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1713335925
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_91
timestamp 1713335925
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_98
timestamp 1713335925
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_114
timestamp 1713335925
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_124
timestamp 1713335925
transform 1 0 12512 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1713335925
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 1713335925
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 1713335925
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 1713335925
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_33
timestamp 1713335925
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_44
timestamp 1713335925
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_62
timestamp 1713335925
transform 1 0 6808 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_74
timestamp 1713335925
transform 1 0 7912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_82
timestamp 1713335925
transform 1 0 8648 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 1713335925
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1713335925
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_120
timestamp 1713335925
transform 1 0 12144 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_136
timestamp 1713335925
transform 1 0 13616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_142
timestamp 1713335925
transform 1 0 14168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 1713335925
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1713335925
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_33
timestamp 1713335925
transform 1 0 4140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_39
timestamp 1713335925
transform 1 0 4692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_47
timestamp 1713335925
transform 1 0 5428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_55
timestamp 1713335925
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_60
timestamp 1713335925
transform 1 0 6624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 1713335925
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 1713335925
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_105
timestamp 1713335925
transform 1 0 10764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_113
timestamp 1713335925
transform 1 0 11500 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_122
timestamp 1713335925
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_134
timestamp 1713335925
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1713335925
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1713335925
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_18
timestamp 1713335925
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_47
timestamp 1713335925
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_57
timestamp 1713335925
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_76
timestamp 1713335925
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_80
timestamp 1713335925
transform 1 0 8464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_88
timestamp 1713335925
transform 1 0 9200 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_92
timestamp 1713335925
transform 1 0 9568 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_100
timestamp 1713335925
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1713335925
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_121
timestamp 1713335925
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_142
timestamp 1713335925
transform 1 0 14168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1713335925
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 1713335925
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_24
timestamp 1713335925
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1713335925
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_41
timestamp 1713335925
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_60
timestamp 1713335925
transform 1 0 6624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1713335925
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_119
timestamp 1713335925
transform 1 0 12052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1713335925
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1713335925
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1713335925
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_6
timestamp 1713335925
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_11
timestamp 1713335925
transform 1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_19
timestamp 1713335925
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_23
timestamp 1713335925
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_27
timestamp 1713335925
transform 1 0 3588 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_29
timestamp 1713335925
transform 1 0 3772 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_35
timestamp 1713335925
transform 1 0 4324 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_43
timestamp 1713335925
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_47
timestamp 1713335925
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1713335925
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_60
timestamp 1713335925
transform 1 0 6624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_71
timestamp 1713335925
transform 1 0 7636 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_79
timestamp 1713335925
transform 1 0 8372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 1713335925
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_85
timestamp 1713335925
transform 1 0 8924 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_91
timestamp 1713335925
transform 1 0 9476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_95
timestamp 1713335925
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_99
timestamp 1713335925
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 1713335925
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1713335925
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_113
timestamp 1713335925
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_119
timestamp 1713335925
transform 1 0 12052 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_127
timestamp 1713335925
transform 1 0 12788 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_131
timestamp 1713335925
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_135
timestamp 1713335925
transform 1 0 13524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_141
timestamp 1713335925
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1713335925
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1713335925
transform 1 0 12880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1713335925
transform -1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1713335925
transform 1 0 11776 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output5
timestamp 1713335925
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1713335925
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1713335925
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1713335925
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1713335925
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 1713335925
transform -1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1713335925
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output12
timestamp 1713335925
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1713335925
transform 1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output14
timestamp 1713335925
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1713335925
transform 1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1713335925
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1713335925
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output18
timestamp 1713335925
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1713335925
transform 1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1713335925
transform 1 0 4048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1713335925
transform 1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output22
timestamp 1713335925
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1713335925
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output24
timestamp 1713335925
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_24
timestamp 1713335925
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1713335925
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_25
timestamp 1713335925
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1713335925
transform -1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_26
timestamp 1713335925
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1713335925
transform -1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_27
timestamp 1713335925
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1713335925
transform -1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_28
timestamp 1713335925
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1713335925
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_29
timestamp 1713335925
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1713335925
transform -1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_30
timestamp 1713335925
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1713335925
transform -1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_31
timestamp 1713335925
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1713335925
transform -1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_32
timestamp 1713335925
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1713335925
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_33
timestamp 1713335925
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1713335925
transform -1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_34
timestamp 1713335925
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1713335925
transform -1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_35
timestamp 1713335925
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1713335925
transform -1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_36
timestamp 1713335925
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1713335925
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_37
timestamp 1713335925
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1713335925
transform -1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_38
timestamp 1713335925
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1713335925
transform -1 0 14536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_39
timestamp 1713335925
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1713335925
transform -1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_40
timestamp 1713335925
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1713335925
transform -1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_41
timestamp 1713335925
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1713335925
transform -1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_42
timestamp 1713335925
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1713335925
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_43
timestamp 1713335925
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1713335925
transform -1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_44
timestamp 1713335925
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1713335925
transform -1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_45
timestamp 1713335925
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1713335925
transform -1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_46
timestamp 1713335925
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1713335925
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_47
timestamp 1713335925
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1713335925
transform -1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 1713335925
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 1713335925
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp 1713335925
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp 1713335925
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp 1713335925
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_53
timestamp 1713335925
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_54
timestamp 1713335925
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp 1713335925
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_56
timestamp 1713335925
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp 1713335925
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp 1713335925
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp 1713335925
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp 1713335925
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp 1713335925
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp 1713335925
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_63
timestamp 1713335925
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_64
timestamp 1713335925
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_65
timestamp 1713335925
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_66
timestamp 1713335925
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp 1713335925
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_68
timestamp 1713335925
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_69
timestamp 1713335925
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_70
timestamp 1713335925
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_71
timestamp 1713335925
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_72
timestamp 1713335925
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_73
timestamp 1713335925
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_74
timestamp 1713335925
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_75
timestamp 1713335925
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_76
timestamp 1713335925
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp 1713335925
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_78
timestamp 1713335925
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_79
timestamp 1713335925
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_80
timestamp 1713335925
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_81
timestamp 1713335925
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_82
timestamp 1713335925
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_83
timestamp 1713335925
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_84
timestamp 1713335925
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_85
timestamp 1713335925
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_86
timestamp 1713335925
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_87
timestamp 1713335925
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_88
timestamp 1713335925
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_89
timestamp 1713335925
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_90
timestamp 1713335925
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_91
timestamp 1713335925
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_92
timestamp 1713335925
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_93
timestamp 1713335925
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_94
timestamp 1713335925
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_95
timestamp 1713335925
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_96
timestamp 1713335925
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_97
timestamp 1713335925
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_98
timestamp 1713335925
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_99
timestamp 1713335925
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_100
timestamp 1713335925
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_101
timestamp 1713335925
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp 1713335925
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_103
timestamp 1713335925
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_104
timestamp 1713335925
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_105
timestamp 1713335925
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_106
timestamp 1713335925
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_107
timestamp 1713335925
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_108
timestamp 1713335925
transform 1 0 3680 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_109
timestamp 1713335925
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_110
timestamp 1713335925
transform 1 0 8832 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_111
timestamp 1713335925
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_112
timestamp 1713335925
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
<< labels >>
rlabel metal1 s 7820 15232 7820 15232 4 VGND
rlabel metal1 s 7820 14688 7820 14688 4 VPWR
rlabel metal2 s 2341 7786 2341 7786 4 _000_
rlabel metal1 s 4181 6698 4181 6698 4 _001_
rlabel metal1 s 6844 13906 6844 13906 4 _002_
rlabel metal1 s 5198 13430 5198 13430 4 _003_
rlabel metal1 s 3854 13974 3854 13974 4 _004_
rlabel metal2 s 2254 14178 2254 14178 4 _005_
rlabel metal2 s 1702 13090 1702 13090 4 _006_
rlabel metal1 s 13008 9554 13008 9554 4 _007_
rlabel metal1 s 9966 8874 9966 8874 4 _008_
rlabel metal1 s 8985 13226 8985 13226 4 _009_
rlabel metal1 s 10794 14314 10794 14314 4 _010_
rlabel metal1 s 12967 10710 12967 10710 4 _011_
rlabel metal1 s 12469 14042 12469 14042 4 _012_
rlabel metal2 s 2438 6120 2438 6120 4 _013_
rlabel metal2 s 2070 4386 2070 4386 4 _014_
rlabel metal2 s 2525 2414 2525 2414 4 _015_
rlabel metal1 s 3629 3026 3629 3026 4 _016_
rlabel metal1 s 4968 2618 4968 2618 4 _017_
rlabel metal2 s 6394 3298 6394 3298 4 _018_
rlabel metal1 s 6036 5202 6036 5202 4 _019_
rlabel metal2 s 7493 2414 7493 2414 4 _020_
rlabel metal1 s 11220 6426 11220 6426 4 _021_
rlabel metal1 s 10610 4522 10610 4522 4 _022_
rlabel metal1 s 6108 6766 6108 6766 4 _023_
rlabel metal1 s 9246 13838 9246 13838 4 _024_
rlabel metal2 s 12829 5678 12829 5678 4 _025_
rlabel metal2 s 12834 4386 12834 4386 4 _026_
rlabel metal1 s 7942 3094 7942 3094 4 _027_
rlabel metal1 s 9414 2346 9414 2346 4 _028_
rlabel metal1 s 8556 14042 8556 14042 4 _029_
rlabel metal2 s 1794 9826 1794 9826 4 _030_
rlabel metal1 s 10863 12206 10863 12206 4 _031_
rlabel metal1 s 6946 8908 6946 8908 4 _032_
rlabel metal1 s 9292 5882 9292 5882 4 _033_
rlabel metal1 s 9154 6698 9154 6698 4 _034_
rlabel metal2 s 6394 7276 6394 7276 4 _035_
rlabel metal1 s 4186 8976 4186 8976 4 _036_
rlabel metal1 s 2622 10744 2622 10744 4 _037_
rlabel metal1 s 6302 7718 6302 7718 4 _038_
rlabel metal1 s 3588 9554 3588 9554 4 _039_
rlabel metal1 s 2346 8874 2346 8874 4 _040_
rlabel metal1 s 2599 9078 2599 9078 4 _041_
rlabel metal1 s 2530 8534 2530 8534 4 _042_
rlabel metal1 s 5888 7854 5888 7854 4 _043_
rlabel metal1 s 6624 8058 6624 8058 4 _044_
rlabel metal1 s 6164 7786 6164 7786 4 _045_
rlabel metal1 s 5415 7922 5415 7922 4 _046_
rlabel metal2 s 3818 7855 3818 7855 4 _047_
rlabel metal1 s 3913 7514 3913 7514 4 _048_
rlabel metal1 s 5750 13910 5750 13910 4 _049_
rlabel metal1 s 6486 9418 6486 9418 4 _050_
rlabel metal1 s 5382 13158 5382 13158 4 _051_
rlabel metal1 s 6026 12138 6026 12138 4 _052_
rlabel metal1 s 5106 11084 5106 11084 4 _053_
rlabel metal1 s 6118 12682 6118 12682 4 _054_
rlabel metal1 s 10580 7378 10580 7378 4 _055_
rlabel metal1 s 10304 7174 10304 7174 4 _056_
rlabel metal1 s 12834 9010 12834 9010 4 _057_
rlabel metal1 s 9752 13906 9752 13906 4 _058_
rlabel metal1 s 6670 12852 6670 12852 4 _059_
rlabel metal1 s 6256 13294 6256 13294 4 _060_
rlabel metal1 s 6210 13702 6210 13702 4 _061_
rlabel metal1 s 2622 11084 2622 11084 4 _062_
rlabel metal1 s 7084 11322 7084 11322 4 _063_
rlabel metal2 s 4922 12653 4922 12653 4 _064_
rlabel metal1 s 5382 13265 5382 13265 4 _065_
rlabel metal1 s 5060 13498 5060 13498 4 _066_
rlabel metal1 s 5612 11118 5612 11118 4 _067_
rlabel metal1 s 5382 10778 5382 10778 4 _068_
rlabel metal1 s 3864 13294 3864 13294 4 _069_
rlabel metal1 s 3726 13498 3726 13498 4 _070_
rlabel metal1 s 4868 11866 4868 11866 4 _071_
rlabel metal1 s 3128 13294 3128 13294 4 _072_
rlabel metal2 s 3174 13600 3174 13600 4 _073_
rlabel metal1 s 11546 9928 11546 9928 4 _074_
rlabel metal1 s 4232 11118 4232 11118 4 _075_
rlabel metal2 s 3174 11764 3174 11764 4 _076_
rlabel metal1 s 2208 12138 2208 12138 4 _077_
rlabel metal1 s 2438 12342 2438 12342 4 _078_
rlabel metal1 s 1794 12818 1794 12818 4 _079_
rlabel metal2 s 9752 11118 9752 11118 4 _080_
rlabel metal1 s 10350 12852 10350 12852 4 _081_
rlabel metal2 s 9982 10489 9982 10489 4 _082_
rlabel metal1 s 12006 9690 12006 9690 4 _083_
rlabel metal1 s 12282 9622 12282 9622 4 _084_
rlabel metal1 s 7038 4012 7038 4012 4 _085_
rlabel metal1 s 9384 13974 9384 13974 4 _086_
rlabel metal1 s 8142 8874 8142 8874 4 _087_
rlabel metal1 s 9246 9010 9246 9010 4 _088_
rlabel metal1 s 10350 10676 10350 10676 4 _089_
rlabel metal1 s 10028 10574 10028 10574 4 _090_
rlabel metal1 s 11362 10506 11362 10506 4 _091_
rlabel metal1 s 11500 10778 11500 10778 4 _092_
rlabel metal1 s 12880 10642 12880 10642 4 _093_
rlabel metal1 s 10258 10608 10258 10608 4 _094_
rlabel metal1 s 9752 10778 9752 10778 4 _095_
rlabel metal2 s 11822 13600 11822 13600 4 _096_
rlabel metal1 s 11040 12750 11040 12750 4 _097_
rlabel metal1 s 10856 12410 10856 12410 4 _098_
rlabel metal1 s 11546 12172 11546 12172 4 _099_
rlabel metal1 s 12650 11628 12650 11628 4 _100_
rlabel metal1 s 11316 13702 11316 13702 4 _101_
rlabel metal2 s 10534 14518 10534 14518 4 _102_
rlabel metal1 s 13662 12138 13662 12138 4 _103_
rlabel metal1 s 12466 11696 12466 11696 4 _104_
rlabel metal2 s 12006 13124 12006 13124 4 _105_
rlabel metal1 s 11822 12274 11822 12274 4 _106_
rlabel metal1 s 12834 12342 12834 12342 4 _107_
rlabel metal1 s 13156 11594 13156 11594 4 _108_
rlabel metal2 s 12282 13940 12282 13940 4 _109_
rlabel metal1 s 12604 14042 12604 14042 4 _110_
rlabel metal1 s 13386 12410 13386 12410 4 _111_
rlabel metal1 s 12696 12954 12696 12954 4 _112_
rlabel metal2 s 7866 5304 7866 5304 4 _113_
rlabel metal1 s 7406 5678 7406 5678 4 _114_
rlabel metal2 s 6578 5406 6578 5406 4 _115_
rlabel metal1 s 6716 4522 6716 4522 4 _116_
rlabel metal1 s 3726 5882 3726 5882 4 _117_
rlabel metal1 s 2691 5678 2691 5678 4 _118_
rlabel metal1 s 3956 5202 3956 5202 4 _119_
rlabel metal2 s 3358 4556 3358 4556 4 _120_
rlabel metal1 s 3634 4114 3634 4114 4 _121_
rlabel metal1 s 3082 3502 3082 3502 4 _122_
rlabel metal1 s 4646 3536 4646 3536 4 _123_
rlabel metal1 s 4094 2414 4094 2414 4 _124_
rlabel metal1 s 5612 4114 5612 4114 4 _125_
rlabel metal1 s 5428 2414 5428 2414 4 _126_
rlabel metal1 s 5750 3604 5750 3604 4 _127_
rlabel metal1 s 6256 3026 6256 3026 4 _128_
rlabel metal1 s 5290 5882 5290 5882 4 _129_
rlabel metal1 s 5796 6290 5796 6290 4 _130_
rlabel metal1 s 7130 4114 7130 4114 4 _131_
rlabel metal1 s 7544 3502 7544 3502 4 _132_
rlabel metal2 s 8418 4590 8418 4590 4 _133_
rlabel metal1 s 10764 5202 10764 5202 4 _134_
rlabel metal1 s 10764 4114 10764 4114 4 _135_
rlabel metal1 s 11546 5644 11546 5644 4 _136_
rlabel metal1 s 9982 5712 9982 5712 4 _137_
rlabel metal1 s 11224 6086 11224 6086 4 _138_
rlabel metal1 s 11454 5814 11454 5814 4 _139_
rlabel metal1 s 9200 5338 9200 5338 4 _140_
rlabel metal1 s 9798 5610 9798 5610 4 _141_
rlabel metal1 s 7084 5882 7084 5882 4 _142_
rlabel metal1 s 12236 5882 12236 5882 4 _143_
rlabel metal1 s 14582 4896 14582 4896 4 _144_
rlabel metal2 s 12282 4760 12282 4760 4 _145_
rlabel metal1 s 12558 4114 12558 4114 4 _146_
rlabel metal2 s 8970 4386 8970 4386 4 _147_
rlabel metal1 s 8786 4454 8786 4454 4 _148_
rlabel metal1 s 9660 3978 9660 3978 4 _149_
rlabel metal1 s 9614 4080 9614 4080 4 _150_
rlabel metal1 s 4324 10778 4324 10778 4 _151_
rlabel metal1 s 2852 10642 2852 10642 4 _152_
rlabel metal1 s 2208 10778 2208 10778 4 _153_
rlabel metal1 s 2162 11254 2162 11254 4 _154_
rlabel metal1 s 1932 9554 1932 9554 4 _155_
rlabel metal1 s 9384 5202 9384 5202 4 _156_
rlabel metal1 s 5980 8262 5980 8262 4 _157_
rlabel metal1 s 2530 13974 2530 13974 4 _158_
rlabel metal1 s 4462 10030 4462 10030 4 _159_
rlabel metal2 s 5764 9554 5764 9554 4 _160_
rlabel metal2 s 8786 12517 8786 12517 4 _161_
rlabel metal1 s 7084 12410 7084 12410 4 _162_
rlabel metal1 s 12926 8398 12926 8398 4 _163_
rlabel metal1 s 5152 9622 5152 9622 4 _164_
rlabel metal1 s 6762 10064 6762 10064 4 _165_
rlabel metal1 s 8832 12410 8832 12410 4 _166_
rlabel metal1 s 9476 7378 9476 7378 4 _167_
rlabel metal1 s 7682 10098 7682 10098 4 _168_
rlabel metal2 s 6946 10336 6946 10336 4 _169_
rlabel metal1 s 6348 10506 6348 10506 4 _170_
rlabel metal2 s 8418 8296 8418 8296 4 _171_
rlabel metal1 s 6670 10608 6670 10608 4 _172_
rlabel metal1 s 4278 9962 4278 9962 4 _173_
rlabel metal1 s 5290 11186 5290 11186 4 _174_
rlabel metal1 s 9936 9622 9936 9622 4 _175_
rlabel metal1 s 5014 12172 5014 12172 4 _176_
rlabel metal1 s 6808 12342 6808 12342 4 _177_
rlabel metal1 s 2714 12104 2714 12104 4 _178_
rlabel metal2 s 3358 9690 3358 9690 4 _179_
rlabel metal1 s 5014 7922 5014 7922 4 _180_
rlabel metal1 s 10902 12138 10902 12138 4 _181_
rlabel metal1 s 6118 7888 6118 7888 4 _182_
rlabel metal1 s 13202 5236 13202 5236 4 _183_
rlabel metal1 s 12052 6290 12052 6290 4 _184_
rlabel metal2 s 12650 8670 12650 8670 4 _185_
rlabel metal1 s 4600 8058 4600 8058 4 _186_
rlabel metal1 s 8372 6358 8372 6358 4 _187_
rlabel metal1 s 7590 6766 7590 6766 4 _188_
rlabel metal1 s 14260 3162 14260 3162 4 adc.comparator.compres.ffsync.stage0
rlabel metal2 s 10902 6018 10902 6018 4 adc.comparator.compres.ffsync.stage1
rlabel metal2 s 13202 9656 13202 9656 4 adc.internalCounter\[0\]
rlabel metal1 s 11040 8942 11040 8942 4 adc.internalCounter\[1\]
rlabel metal1 s 7544 12206 7544 12206 4 adc.internalCounter\[2\]
rlabel metal1 s 11730 13940 11730 13940 4 adc.internalCounter\[3\]
rlabel metal1 s 13938 12240 13938 12240 4 adc.internalCounter\[4\]
rlabel metal1 s 13708 12954 13708 12954 4 adc.internalCounter\[5\]
rlabel metal1 s 11454 6868 11454 6868 4 adc.state\[0\]
rlabel metal2 s 9614 7378 9614 7378 4 adc.state\[1\]
rlabel metal1 s 8280 7174 8280 7174 4 adc.state\[2\]
rlabel metal2 s 10442 13333 10442 13333 4 adc.state\[3\]
rlabel metal1 s 9108 3162 9108 3162 4 adc.syncroCount\[0\]
rlabel metal1 s 10580 2618 10580 2618 4 adc.syncroCount\[1\]
rlabel metal2 s 14950 1554 14950 1554 4 analog_comparator_out
rlabel metal1 s 12880 14994 12880 14994 4 calib_enable
rlabel metal2 s 15042 12845 15042 12845 4 clk
rlabel metal1 s 7360 8398 7360 8398 4 clknet_0_clk
rlabel metal1 s 1978 2482 1978 2482 4 clknet_2_0__leaf_clk
rlabel metal1 s 1794 7922 1794 7922 4 clknet_2_1__leaf_clk
rlabel metal1 s 9798 2414 9798 2414 4 clknet_2_2__leaf_clk
rlabel metal1 s 12558 10506 12558 10506 4 clknet_2_3__leaf_clk
rlabel metal2 s 13662 959 13662 959 4 comparator_nen
rlabel metal2 s 782 1520 782 1520 4 dac_set[0]
rlabel metal2 s 2070 1520 2070 1520 4 dac_set[1]
rlabel metal2 s 3358 823 3358 823 4 dac_set[2]
rlabel metal2 s 4646 1520 4646 1520 4 dac_set[3]
rlabel metal2 s 5934 1520 5934 1520 4 dac_set[4]
rlabel metal2 s 7222 959 7222 959 4 dac_set[5]
rlabel metal2 s 8510 959 8510 959 4 dac_set[6]
rlabel metal2 s 9798 1554 9798 1554 4 dac_set[7]
rlabel metal2 s 12374 1520 12374 1520 4 do_calibrate
rlabel metal1 s 13197 3026 13197 3026 4 net1
rlabel metal1 s 6118 2414 6118 2414 4 net10
rlabel metal1 s 7176 3366 7176 3366 4 net11
rlabel metal1 s 8970 2414 8970 2414 4 net12
rlabel metal1 s 10672 2414 10672 2414 4 net13
rlabel metal1 s 13524 2482 13524 2482 4 net14
rlabel metal1 s 7958 14042 7958 14042 4 net15
rlabel metal1 s 4646 13906 4646 13906 4 net16
rlabel metal1 s 4876 14042 4876 14042 4 net17
rlabel metal2 s 3266 14722 3266 14722 4 net18
rlabel metal1 s 2806 13260 2806 13260 4 net19
rlabel metal2 s 13202 14790 13202 14790 4 net2
rlabel metal2 s 4278 13707 4278 13707 4 net20
rlabel metal1 s 3312 14994 3312 14994 4 net21
rlabel metal1 s 2070 15028 2070 15028 4 net22
rlabel metal2 s 1610 14790 1610 14790 4 net23
rlabel metal1 s 11224 2414 11224 2414 4 net24
rlabel metal2 s 2990 8738 2990 8738 4 net3
rlabel metal2 s 13570 4862 13570 4862 4 net4
rlabel metal1 s 14214 2414 14214 2414 4 net5
rlabel metal1 s 2484 6086 2484 6086 4 net6
rlabel metal1 s 2254 2414 2254 2414 4 net7
rlabel metal1 s 4324 2414 4324 2414 4 net8
rlabel metal1 s 4738 2414 4738 2414 4 net9
rlabel metal1 s 9568 15130 9568 15130 4 result[0]
rlabel metal2 s 8510 16167 8510 16167 4 result[1]
rlabel metal2 s 7406 16167 7406 16167 4 result[2]
rlabel metal1 s 6302 15130 6302 15130 4 result[3]
rlabel metal1 s 5290 15130 5290 15130 4 result[4]
rlabel metal1 s 4048 15130 4048 15130 4 result[5]
rlabel metal1 s 2944 15130 2944 15130 4 result[6]
rlabel metal2 s 1886 16167 1886 16167 4 result[7]
rlabel metal1 s 1058 15130 1058 15130 4 result_ready
rlabel metal2 s 13938 16092 13938 16092 4 rst
rlabel metal2 s 11086 823 11086 823 4 thresh_sel
rlabel metal4 s 10603 13668 10603 13668 4 use_ext_thresh
rlabel metal1 s 11776 14994 11776 14994 4 user_enable
flabel metal4 s 10904 2128 11304 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4904 2128 5304 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13904 2128 14304 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7904 2128 8304 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1904 2128 2304 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 14922 0 14978 800 0 FreeSans 280 90 0 0 analog_comparator_out
port 3 nsew
flabel metal2 s 12806 17064 12862 17864 0 FreeSans 280 90 0 0 calib_enable
port 4 nsew
flabel metal2 s 15014 17064 15070 17864 0 FreeSans 280 90 0 0 clk
port 5 nsew
flabel metal2 s 13634 0 13690 800 0 FreeSans 280 90 0 0 comparator_nen
port 6 nsew
flabel metal2 s 754 0 810 800 0 FreeSans 280 90 0 0 dac_set[0]
port 7 nsew
flabel metal2 s 2042 0 2098 800 0 FreeSans 280 90 0 0 dac_set[1]
port 8 nsew
flabel metal2 s 3330 0 3386 800 0 FreeSans 280 90 0 0 dac_set[2]
port 9 nsew
flabel metal2 s 4618 0 4674 800 0 FreeSans 280 90 0 0 dac_set[3]
port 10 nsew
flabel metal2 s 5906 0 5962 800 0 FreeSans 280 90 0 0 dac_set[4]
port 11 nsew
flabel metal2 s 7194 0 7250 800 0 FreeSans 280 90 0 0 dac_set[5]
port 12 nsew
flabel metal2 s 8482 0 8538 800 0 FreeSans 280 90 0 0 dac_set[6]
port 13 nsew
flabel metal2 s 9770 0 9826 800 0 FreeSans 280 90 0 0 dac_set[7]
port 14 nsew
flabel metal2 s 12346 0 12402 800 0 FreeSans 280 90 0 0 do_calibrate
port 15 nsew
flabel metal2 s 9494 17064 9550 17864 0 FreeSans 280 90 0 0 result[0]
port 16 nsew
flabel metal2 s 8390 17064 8446 17864 0 FreeSans 280 90 0 0 result[1]
port 17 nsew
flabel metal2 s 7286 17064 7342 17864 0 FreeSans 280 90 0 0 result[2]
port 18 nsew
flabel metal2 s 6182 17064 6238 17864 0 FreeSans 280 90 0 0 result[3]
port 19 nsew
flabel metal2 s 5078 17064 5134 17864 0 FreeSans 280 90 0 0 result[4]
port 20 nsew
flabel metal2 s 3974 17064 4030 17864 0 FreeSans 280 90 0 0 result[5]
port 21 nsew
flabel metal2 s 2870 17064 2926 17864 0 FreeSans 280 90 0 0 result[6]
port 22 nsew
flabel metal2 s 1766 17064 1822 17864 0 FreeSans 280 90 0 0 result[7]
port 23 nsew
flabel metal2 s 662 17064 718 17864 0 FreeSans 280 90 0 0 result_ready
port 24 nsew
flabel metal2 s 13910 17064 13966 17864 0 FreeSans 280 90 0 0 rst
port 25 nsew
flabel metal2 s 11058 0 11114 800 0 FreeSans 280 90 0 0 thresh_sel
port 26 nsew
flabel metal2 s 10598 17064 10654 17864 0 FreeSans 280 90 0 0 use_ext_thresh
port 27 nsew
flabel metal2 s 11702 17064 11758 17864 0 FreeSans 280 90 0 0 user_enable
port 28 nsew
<< properties >>
string FIXED_BBOX 0 0 15720 17864
string GDS_END 1119870
string GDS_FILE wowa_digital_ol.gds
string GDS_START 439436
<< end >>
