magic
tech sky130A
magscale 1 2
timestamp 1713420955
<< metal1 >>
rect 5630 5350 6440 5620
rect 5630 4575 5900 5350
rect 6074 5164 6332 5256
rect 6074 4290 6166 5164
rect 6200 4520 6400 4720
rect 7000 4520 7200 4720
rect 5240 4090 5440 4290
rect 5840 4094 6166 4290
rect 5840 4090 6150 4094
rect 6140 3977 6240 4020
rect 6125 3858 6131 3977
rect 6250 3858 6357 3977
rect 6140 3820 6240 3858
rect 5240 3520 6400 3740
<< via1 >>
rect 6131 3858 6250 3977
<< metal2 >>
rect 5745 4290 6266 4295
rect 5240 4144 6266 4290
rect 5240 4090 5960 4144
rect 6115 3977 6266 4144
rect 6115 3858 6131 3977
rect 6250 3858 6266 3977
rect 6115 3842 6266 3858
use lvtnot  x1
timestamp 1713420648
transform 1 0 3820 0 1 3390
box 1400 340 2238 1340
use passgate  x2
timestamp 1713420955
transform 1 0 4000 0 1 4220
box 2200 -700 3200 1400
<< labels >>
flabel metal1 6200 4520 6400 4720 0 FreeSans 1280 0 0 0 IN
port 1 nsew
flabel metal1 7000 4520 7200 4720 0 FreeSans 1280 0 0 0 OUT
port 2 nsew
flabel metal1 5240 4090 5440 4290 0 FreeSans 1280 0 0 0 EN
port 0 nsew
flabel metal1 5910 5360 6110 5560 0 FreeSans 1280 0 0 0 VCC
port 3 nsew
flabel metal1 5910 3520 6110 3720 0 FreeSans 1280 0 0 0 VSS
port 4 nsew
<< end >>
