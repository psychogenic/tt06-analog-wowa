magic
tech sky130A
magscale 1 2
timestamp 1713420648
<< pwell >>
rect 1740 560 1880 600
rect 1710 550 1880 560
rect 1680 500 1880 550
rect 1680 480 1740 500
<< locali >>
rect 1420 460 1560 670
rect 1420 430 1620 460
rect 2070 460 2160 670
rect 2010 430 2160 460
rect 1420 340 2160 430
<< viali >>
rect 1620 1220 2010 1270
rect 1620 430 2010 480
<< metal1 >>
rect 1420 1270 2160 1340
rect 1420 1220 1620 1270
rect 2010 1220 2160 1270
rect 1420 1140 2160 1220
rect 1520 1100 1580 1110
rect 2060 1100 2120 1110
rect 1500 1040 1510 1100
rect 1580 1040 1590 1100
rect 2050 1040 2060 1100
rect 2130 1040 2140 1100
rect 1520 1030 1580 1040
rect 2060 1030 2120 1040
rect 1420 885 1620 900
rect 1420 715 1430 885
rect 1600 715 1620 885
rect 1420 700 1620 715
rect 1730 880 1880 1030
rect 2020 880 2220 900
rect 1730 750 2220 880
rect 1620 640 1680 650
rect 1590 580 1600 640
rect 1670 580 1680 640
rect 1730 630 1880 750
rect 2020 700 2220 750
rect 1950 640 2010 660
rect 1740 580 1880 600
rect 1940 580 1950 640
rect 2020 580 2030 640
rect 1720 560 1900 580
rect 1710 550 1900 560
rect 1420 520 1620 540
rect 1680 520 1940 550
rect 1420 480 2160 520
rect 1420 430 1620 480
rect 2010 430 2160 480
rect 1420 340 2160 430
<< via1 >>
rect 1510 1040 1580 1100
rect 2060 1040 2130 1100
rect 1430 715 1600 885
rect 1600 580 1670 640
rect 1950 580 2020 640
<< metal2 >>
rect 1430 1100 2160 1130
rect 1430 1040 1510 1100
rect 1580 1040 2060 1100
rect 2130 1040 2160 1100
rect 1430 1010 2160 1040
rect 1430 885 1600 1010
rect 1430 670 1600 715
rect 1430 640 2160 670
rect 1430 580 1600 640
rect 1670 580 1950 640
rect 2020 580 2160 640
rect 1430 550 2160 580
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1
timestamp 1713125502
transform 0 -1 1810 1 0 611
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QFWD3  XM2
timestamp 1713125502
transform 0 1 1819 -1 0 1071
box -231 -419 231 419
<< labels >>
flabel metal1 1420 700 1620 900 0 FreeSans 1280 0 0 0 a
port 0 nsew
flabel metal1 2020 700 2220 900 0 FreeSans 1280 0 0 0 y
port 1 nsew
flabel metal1 1420 1140 1620 1340 0 FreeSans 1280 0 0 0 VCCPIN
port 2 nsew
flabel metal1 1420 340 1620 540 0 FreeSans 1280 0 0 0 VSSPIN
port 3 nsew
<< end >>
