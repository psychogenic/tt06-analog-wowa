* NGSPICE file created from wowa_analog_parax.ext - technology: sky130A

.subckt wowa_analog_parax b0 b1 b2 b3 b4 b5 b6 b7 EXTTHRESH USEEXT DACOUT INPUT VCC
+ CAL VSS COMPOUT EN_N
X0 a_6766_30798# a_7366_26366# VSS.t4 sky130_fd_pr__res_high_po_0p35 l=20.16
X1 x1.x1.pg2g.t1 x1.x1.pg2g.t0 x1.x1.mirhigh.t1 VCC.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
X2 x1.x2.OUT.t1 x1.x2.x2.GP COMPOUT.t2 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X3 a_5366_34798# VSS VSS.t32 sky130_fd_pr__res_high_po_0p35 l=40.16
X4 x1.x2.OUT.t0 CAL.t0 COMPOUT.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X5 x1.x3.SEL_N.t1 CAL.t1 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6 VCC.t19 EN_N.t0 x1.x1.mirhigh.t2 VCC.t18 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.15
X7 x1.x1.G2 x1.x1.G2 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X8 a_9166_30798# a_8566_26366# VSS.t6 sky130_fd_pr__res_high_po_0p35 l=20.16
X9 x3.SEL_N.t0 USEEXT.t0 VCC.t10 VCC.t9 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
X10 b2 a_6766_30798# VSS.t4 sky130_fd_pr__res_high_po_0p35 l=40.16
X11 VSS.t31 x1.x1.G1 x1.x1.G1 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X12 x1.x2.OUT.t2 VSS.t13 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X13 a_5366_34798# a_6166_26366# VSS.t16 sky130_fd_pr__res_high_po_0p35 l=20.16
X14 x3.OUT.t5 x1.x3.SEL_N.t2 x1.x3.OUT.t2 VCC.t14 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X15 x1.x1.n2n VCC.t22 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X16 x1.x1.G2 x1.x3.OUT.t4 x1.x1.inhigh.t1 VCC.t15 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
X17 b5 a_8566_26366# VSS.t6 sky130_fd_pr__res_high_po_0p35 l=40.16
X18 b7 DACOUT VSS.t38 sky130_fd_pr__res_high_po_0p35 l=40.16
X19 VCC.t12 EN_N.t1 x1.x1.p2p VCC.t11 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X20 VSS.t23 EN_N.t2 COMPOUT.t3 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X21 x3.OUT.t2 x3.SEL_N.t2 EXTTHRESH.t0 VCC.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X22 x1.x2.x2.Z VSS.t15 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X23 b0 a_5366_34798# VSS.t16 sky130_fd_pr__res_high_po_0p35 l=40.16
X24 x1.x1.inhigh.t0 x3.OUT.t6 x1.x1.G1 VCC.t21 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
X25 VCC.t8 CAL.t2 x1.x2.x2.GP VCC.t7 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
X26 a_7966_30798# a_7366_26366# VSS.t11 sky130_fd_pr__res_high_po_0p35 l=20.16
X27 x1.x2.x2.Z VSS.t14 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X28 x3.OUT.t4 USEEXT.t1 EXTTHRESH.t1 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X29 x1.x2.x2.GP CAL.t3 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X30 a_9166_30798# DACOUT VSS.t8 sky130_fd_pr__res_high_po_0p35 l=20.16
X31 b3 a_7366_26366# VSS.t11 sky130_fd_pr__res_high_po_0p35 l=40.16
X32 a_6766_30798# a_6166_26366# VSS.t7 sky130_fd_pr__res_high_po_0p35 l=20.16
X33 x1.x1.mirhigh.t0 x1.x1.pg2g.t2 COMPOUT.t4 VCC.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
X34 x1.x1.pg2g x1.x1.G1 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X35 x3.OUT.t1 x3.SEL_N.t3 DACOUT.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X36 VCC.t1 CAL.t4 x1.x3.SEL_N.t0 VCC.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
X37 b6 a_9166_30798# VSS.t8 sky130_fd_pr__res_high_po_0p35 l=40.16
X38 VSS.t1 x1.x1.G2 COMPOUT.t0 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X39 x1.x1.inhigh.t2 EN_N.t3 VCC.t3 VCC.t2 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=8
X40 x1.x1.G1 x1.x2.OUT.t3 x1.x1.n2n VSS.t37 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X41 x1.x3.OUT.t3 x1.x3.SEL_N.t3 INPUT.t1 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X42 a_7966_30798# a_8566_26366# VSS.t10 sky130_fd_pr__res_high_po_0p35 l=20.16
X43 VSS.t21 USEEXT.t2 x3.SEL_N.t1 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X44 b1 a_6166_26366# VSS.t7 sky130_fd_pr__res_high_po_0p35 l=40.16
X45 x1.x2.OUT.t2 VSS.t12 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X46 x3.OUT.t0 CAL.t5 x1.x3.OUT.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X47 x3.OUT.t3 USEEXT.t3 DACOUT.t2 VCC.t6 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
X48 b4 a_7966_30798# VSS.t10 sky130_fd_pr__res_high_po_0p35 l=40.16
X49 x1.x1.G1 x1.x2.OUT.t4 x1.x1.p2p VCC.t13 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X50 x1.x3.OUT.t1 CAL.t6 INPUT.t0 VCC.t20 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
R0 VSS.n330 VSS.n156 1.1352e+06
R1 VSS.n302 VSS.n301 88402
R2 VSS.n331 VSS.n330 85360
R3 VSS.n301 VSS.n153 57710.7
R4 VSS.n301 VSS.n293 42701
R5 VSS.n290 VSS.n289 38439
R6 VSS.n417 VSS.n90 37991.8
R7 VSS.n290 VSS.n154 30084.4
R8 VSS.n486 VSS.n3 27093.3
R9 VSS.n8 VSS.n4 27093.3
R10 VSS.n8 VSS.n3 27093.3
R11 VSS.n468 VSS.n27 27093.3
R12 VSS.n468 VSS.n467 27093.3
R13 VSS.n467 VSS.n463 27093.3
R14 VSS.n463 VSS.n27 27093.3
R15 VSS.n472 VSS.n21 27093.3
R16 VSS.n472 VSS.n22 27093.3
R17 VSS.n21 VSS.n20 27093.3
R18 VSS.n22 VSS.n20 27093.3
R19 VSS.n453 VSS.n42 27093.3
R20 VSS.n453 VSS.n43 27093.3
R21 VSS.n42 VSS.n41 27093.3
R22 VSS.n43 VSS.n41 27093.3
R23 VSS.n449 VSS.n46 27093.3
R24 VSS.n449 VSS.n47 27093.3
R25 VSS.n448 VSS.n46 27093.3
R26 VSS.n448 VSS.n47 27093.3
R27 VSS.n437 VSS.n57 27093.3
R28 VSS.n437 VSS.n58 27093.3
R29 VSS.n438 VSS.n57 27093.3
R30 VSS.n438 VSS.n58 27093.3
R31 VSS.n432 VSS.n68 27093.3
R32 VSS.n432 VSS.n69 27093.3
R33 VSS.n431 VSS.n68 27093.3
R34 VSS.n431 VSS.n69 27093.3
R35 VSS.n426 VSS.n78 27093.3
R36 VSS.n426 VSS.n79 27093.3
R37 VSS.n427 VSS.n78 27093.3
R38 VSS.n427 VSS.n79 27093.3
R39 VSS.n422 VSS.n88 27093.3
R40 VSS.n422 VSS.n89 27093.3
R41 VSS.n421 VSS.n88 27093.3
R42 VSS.n421 VSS.n89 27093.3
R43 VSS.n331 VSS.n153 23925
R44 VSS.n326 VSS.n325 20589.7
R45 VSS.n325 VSS.n324 19594.2
R46 VSS.n100 VSS.n99 18357.1
R47 VSS.n301 VSS.n155 17328.1
R48 VSS.n30 VSS.n6 15505.1
R49 VSS.n30 VSS.n7 15505.1
R50 VSS.n483 VSS.n6 15505.1
R51 VSS.n483 VSS.n7 15505.1
R52 VSS.n16 VSS.n13 15505.1
R53 VSS.n16 VSS.n14 15505.1
R54 VSS.n473 VSS.n13 15505.1
R55 VSS.n473 VSS.n14 15505.1
R56 VSS.n454 VSS.n34 15505.1
R57 VSS.n454 VSS.n35 15505.1
R58 VSS.n39 VSS.n34 15505.1
R59 VSS.n39 VSS.n35 15505.1
R60 VSS.n370 VSS.n48 15505.1
R61 VSS.n375 VSS.n48 15505.1
R62 VSS.n370 VSS.n51 15505.1
R63 VSS.n375 VSS.n51 15505.1
R64 VSS.n385 VSS.n60 15505.1
R65 VSS.n368 VSS.n60 15505.1
R66 VSS.n385 VSS.n64 15505.1
R67 VSS.n368 VSS.n64 15505.1
R68 VSS.n392 VSS.n71 15505.1
R69 VSS.n366 VSS.n71 15505.1
R70 VSS.n392 VSS.n74 15505.1
R71 VSS.n366 VSS.n74 15505.1
R72 VSS.n362 VSS.n81 15505.1
R73 VSS.n391 VSS.n81 15505.1
R74 VSS.n362 VSS.n84 15505.1
R75 VSS.n391 VSS.n84 15505.1
R76 VSS.n173 VSS.n163 15252.3
R77 VSS.n163 VSS.n155 14240.6
R78 VSS.n352 VSS.n136 13926.5
R79 VSS.n330 VSS.n155 13892
R80 VSS.n407 VSS.n98 13166.6
R81 VSS.n407 VSS.n90 11573.8
R82 VSS.n325 VSS.n162 10139.7
R83 VSS.n407 VSS.n99 9491.27
R84 VSS.n331 VSS.n154 9075
R85 VSS.n329 VSS.n328 8450.84
R86 VSS.n328 VSS.n98 8440.71
R87 VSS.n327 VSS.n326 7196.9
R88 VSS.n145 VSS.n144 6564.74
R89 VSS.n344 VSS.n144 6564.74
R90 VSS.n344 VSS.n342 6564.74
R91 VSS.n342 VSS.n145 6564.74
R92 VSS.n328 VSS.n327 6540.44
R93 VSS.n327 VSS.n162 5785.42
R94 VSS.n303 VSS.n151 5116.21
R95 VSS.n303 VSS.n152 5116.21
R96 VSS.n333 VSS.n152 5116.21
R97 VSS.n333 VSS.n151 5116.21
R98 VSS.n307 VSS.n178 5116.21
R99 VSS.n307 VSS.n179 5116.21
R100 VSS.n308 VSS.n178 5116.21
R101 VSS.n308 VSS.n179 5116.21
R102 VSS.n322 VSS.n166 5116.21
R103 VSS.n174 VSS.n166 5116.21
R104 VSS.n174 VSS.n167 5116.21
R105 VSS.n322 VSS.n167 5116.21
R106 VSS.n203 VSS.n199 5116.21
R107 VSS.n199 VSS.n169 5116.21
R108 VSS.n200 VSS.n169 5116.21
R109 VSS.n203 VSS.n200 5116.21
R110 VSS.n231 VSS.n156 3851.76
R111 VSS.n180 VSS.n162 3531.49
R112 VSS.n229 VSS.n134 2914.44
R113 VSS.n354 VSS.n134 2914.44
R114 VSS.n229 VSS.n135 2914.44
R115 VSS.n354 VSS.n135 2914.44
R116 VSS.n247 VSS.n227 2914.44
R117 VSS.n256 VSS.n227 2914.44
R118 VSS.n247 VSS.n228 2914.44
R119 VSS.n256 VSS.n228 2914.44
R120 VSS.n287 VSS.n182 2914.44
R121 VSS.n287 VSS.n183 2914.44
R122 VSS.n272 VSS.n182 2914.44
R123 VSS.n272 VSS.n183 2914.44
R124 VSS.n116 VSS.n109 2914.44
R125 VSS.n113 VSS.n109 2914.44
R126 VSS.n113 VSS.n110 2914.44
R127 VSS.n116 VSS.n110 2914.44
R128 VSS.n111 VSS.n101 2914.44
R129 VSS.n405 VSS.n101 2914.44
R130 VSS.n405 VSS.n102 2914.44
R131 VSS.n111 VSS.n102 2914.44
R132 VSS.n157 VSS.n137 2508.85
R133 VSS.n350 VSS.n137 2508.85
R134 VSS.n157 VSS.n138 2508.85
R135 VSS.n350 VSS.n138 2508.85
R136 VSS.n326 VSS.n163 2472.45
R137 VSS.n409 VSS.n91 2306.06
R138 VSS.n415 VSS.n91 2306.06
R139 VSS.n409 VSS.n92 2306.06
R140 VSS.n415 VSS.n92 2306.06
R141 VSS.n244 VSS.n232 2306.06
R142 VSS.n253 VSS.n232 2306.06
R143 VSS.n244 VSS.n233 2306.06
R144 VSS.n253 VSS.n233 2306.06
R145 VSS.n277 VSS.n270 2306.06
R146 VSS.n277 VSS.n271 2306.06
R147 VSS.n278 VSS.n270 2306.06
R148 VSS.n278 VSS.n271 2306.06
R149 VSS.n207 VSS.n195 2306.06
R150 VSS.n208 VSS.n195 2306.06
R151 VSS.n208 VSS.n194 2306.06
R152 VSS.n207 VSS.n194 2306.06
R153 VSS.t0 VSS.n164 2152.43
R154 VSS.n173 VSS.t28 2152.43
R155 VSS.n302 VSS.t30 1874.46
R156 VSS.n332 VSS.t30 1863.35
R157 VSS.n420 VSS.n87 1760.38
R158 VSS.n423 VSS.n87 1760.38
R159 VSS.n201 VSS.n165 1590
R160 VSS.n90 VSS.n83 1477.58
R161 VSS.n196 VSS.n180 1382.33
R162 VSS.n332 VSS.n331 1315.3
R163 VSS.n291 VSS.n290 1306.25
R164 VSS.n160 VSS.n156 1273.43
R165 VSS.t28 VSS.n165 1256.58
R166 VSS.n136 VSS.n98 1052.91
R167 VSS.n289 VSS.n180 910.42
R168 VSS.n323 VSS.n165 895.856
R169 VSS.n351 VSS.n350 823.056
R170 VSS.n324 VSS.n164 761.082
R171 VSS.t2 VSS.n291 678.75
R172 VSS.t32 VSS.n484 647
R173 VSS.n324 VSS.n323 642.163
R174 VSS.t2 VSS.n293 623.75
R175 VSS.n418 VSS.n417 535.436
R176 VSS.n202 VSS.n197 514.71
R177 VSS.n306 VSS.n177 451.89
R178 VSS.n274 VSS.n273 431.83
R179 VSS.n202 VSS.n201 427.839
R180 VSS.n146 VSS.n142 426.541
R181 VSS.n304 VSS.n300 426.505
R182 VSS.n345 VSS.n142 359.279
R183 VSS.n487 VSS.n2 348.882
R184 VSS.n343 VSS.t25 343.591
R185 VSS.n175 VSS.n172 322.786
R186 VSS.n330 VSS.t30 313.719
R187 VSS.n288 VSS.n181 305.168
R188 VSS.n85 VSS.n73 301.67
R189 VSS.n75 VSS.n63 301.67
R190 VSS.n369 VSS.n65 301.67
R191 VSS.n52 VSS.n38 301.67
R192 VSS.n40 VSS.n18 301.67
R193 VSS.n29 VSS.n19 301.67
R194 VSS.n488 VSS.n487 295.498
R195 VSS.n207 VSS.n206 292.5
R196 VSS.t22 VSS.n207 292.5
R197 VSS.n209 VSS.n208 292.5
R198 VSS.n208 VSS.t22 292.5
R199 VSS.n109 VSS.n108 292.5
R200 VSS.t27 VSS.n109 292.5
R201 VSS.n111 VSS.n104 292.5
R202 VSS.n112 VSS.n111 292.5
R203 VSS.n110 VSS.n107 292.5
R204 VSS.t27 VSS.n110 292.5
R205 VSS.n271 VSS.n269 292.5
R206 VSS.n275 VSS.n271 292.5
R207 VSS.n270 VSS.n268 292.5
R208 VSS.n274 VSS.n270 292.5
R209 VSS.n272 VSS.n185 292.5
R210 VSS.t5 VSS.n272 292.5
R211 VSS.n287 VSS.n286 292.5
R212 VSS.n288 VSS.n287 292.5
R213 VSS.n257 VSS.n256 292.5
R214 VSS.n256 VSS.n255 292.5
R215 VSS.n248 VSS.n247 292.5
R216 VSS.n247 VSS.n246 292.5
R217 VSS.n253 VSS.n252 292.5
R218 VSS.n254 VSS.n253 292.5
R219 VSS.n244 VSS.n243 292.5
R220 VSS.n245 VSS.n244 292.5
R221 VSS.n135 VSS.n132 292.5
R222 VSS.t9 VSS.n135 292.5
R223 VSS.n134 VSS.n133 292.5
R224 VSS.t9 VSS.n134 292.5
R225 VSS.n405 VSS.n404 292.5
R226 VSS.n406 VSS.n405 292.5
R227 VSS.n413 VSS.n92 292.5
R228 VSS.n92 VSS.t20 292.5
R229 VSS.n93 VSS.n91 292.5
R230 VSS.n91 VSS.t20 292.5
R231 VSS.n383 VSS.n74 292.5
R232 VSS.t6 VSS.n74 292.5
R233 VSS.n367 VSS.n64 292.5
R234 VSS.t10 VSS.n64 292.5
R235 VSS.n378 VSS.n51 292.5
R236 VSS.t11 VSS.n51 292.5
R237 VSS.n373 VSS.n39 292.5
R238 VSS.t4 VSS.n39 292.5
R239 VSS.n474 VSS.n473 292.5
R240 VSS.n473 VSS.t7 292.5
R241 VSS.n479 VSS.n7 292.5
R242 VSS.n7 VSS.t16 292.5
R243 VSS.n395 VSS.n84 292.5
R244 VSS.t8 VSS.n84 292.5
R245 VSS.n365 VSS.n81 292.5
R246 VSS.t8 VSS.n81 292.5
R247 VSS.n389 VSS.n71 292.5
R248 VSS.t6 VSS.n71 292.5
R249 VSS.n387 VSS.n60 292.5
R250 VSS.t10 VSS.n60 292.5
R251 VSS.n54 VSS.n48 292.5
R252 VSS.t11 VSS.n48 292.5
R253 VSS.n455 VSS.n454 292.5
R254 VSS.n454 VSS.t4 292.5
R255 VSS.n457 VSS.n16 292.5
R256 VSS.t7 VSS.n16 292.5
R257 VSS.n459 VSS.n6 292.5
R258 VSS.n6 VSS.t16 292.5
R259 VSS.n428 VSS.n427 292.5
R260 VSS.n427 VSS.t8 292.5
R261 VSS.n431 VSS.n430 292.5
R262 VSS.t6 VSS.n431 292.5
R263 VSS.n439 VSS.n438 292.5
R264 VSS.n438 VSS.t10 292.5
R265 VSS.n448 VSS.n447 292.5
R266 VSS.t11 VSS.n448 292.5
R267 VSS.n445 VSS.n41 292.5
R268 VSS.t4 VSS.n41 292.5
R269 VSS.n443 VSS.n20 292.5
R270 VSS.t7 VSS.n20 292.5
R271 VSS.n463 VSS.n462 292.5
R272 VSS.n463 VSS.t16 292.5
R273 VSS.n421 VSS.n420 292.5
R274 VSS.t38 VSS.n421 292.5
R275 VSS.n423 VSS.n422 292.5
R276 VSS.n422 VSS.t38 292.5
R277 VSS.n426 VSS.n425 292.5
R278 VSS.t8 VSS.n426 292.5
R279 VSS.n433 VSS.n432 292.5
R280 VSS.n432 VSS.t6 292.5
R281 VSS.n437 VSS.n436 292.5
R282 VSS.t10 VSS.n437 292.5
R283 VSS.n450 VSS.n449 292.5
R284 VSS.n449 VSS.t11 292.5
R285 VSS.n453 VSS.n452 292.5
R286 VSS.t4 VSS.n453 292.5
R287 VSS.n472 VSS.n471 292.5
R288 VSS.t7 VSS.n472 292.5
R289 VSS.n469 VSS.n468 292.5
R290 VSS.n468 VSS.t16 292.5
R291 VSS.n464 VSS.n3 292.5
R292 VSS.t32 VSS.n3 292.5
R293 VSS.n480 VSS.n4 292.5
R294 VSS.n485 VSS.n4 288.712
R295 VSS.n231 VSS.n230 287.026
R296 VSS.n275 VSS.n154 260.13
R297 VSS.n136 VSS.n99 259.06
R298 VSS.n316 VSS.n315 258.839
R299 VSS.n305 VSS.n304 249.601
R300 VSS.n306 VSS.n305 249.601
R301 VSS.n343 VSS.n136 249.587
R302 VSS.n334 VSS.n150 244.138
R303 VSS.n158 VSS.t37 241.245
R304 VSS.n480 VSS.n2 232.353
R305 VSS.n346 VSS.t26 229.185
R306 VSS.n205 VSS.n198 217.103
R307 VSS.n466 VSS.n5 199.749
R308 VSS.n198 VSS.n168 198.024
R309 VSS.n172 VSS.n168 198.024
R310 VSS.n286 VSS.n184 189.365
R311 VSS.n286 VSS.n285 189.365
R312 VSS.n114 VSS.n100 174.674
R313 VSS.t22 VSS.n196 171.571
R314 VSS.t22 VSS.n197 171.571
R315 VSS.n470 VSS.n24 171.476
R316 VSS.n28 VSS.n24 171.476
R317 VSS.n442 VSS.n23 171.476
R318 VSS.n444 VSS.n442 171.476
R319 VSS.n451 VSS.n44 171.476
R320 VSS.n446 VSS.n44 171.476
R321 VSS.n55 VSS.n45 171.476
R322 VSS.n440 VSS.n55 171.476
R323 VSS.n434 VSS.n66 171.476
R324 VSS.n66 VSS.n56 171.476
R325 VSS.n76 VSS.n67 171.476
R326 VSS.n429 VSS.n76 171.476
R327 VSS.n424 VSS.n86 171.476
R328 VSS.n86 VSS.n77 171.476
R329 VSS.t18 VSS.n274 166.637
R330 VSS.t18 VSS.n275 166.637
R331 VSS.n349 VSS.n139 163.012
R332 VSS.n140 VSS.n139 163.012
R333 VSS.n182 VSS.n181 162.441
R334 VSS.n159 VSS.n158 158.845
R335 VSS.n349 VSS.n348 158.72
R336 VSS.n115 VSS.t27 157.766
R337 VSS.n347 VSS.n140 156.988
R338 VSS.n330 VSS.n329 156.124
R339 VSS.t27 VSS.t17 150.99
R340 VSS.n352 VSS.t37 149.911
R341 VSS.t8 VSS.n83 146.865
R342 VSS.t8 VSS.n85 146.865
R343 VSS.t6 VSS.n73 146.865
R344 VSS.t6 VSS.n75 146.865
R345 VSS.t10 VSS.n63 146.865
R346 VSS.t10 VSS.n65 146.865
R347 VSS.t11 VSS.n52 146.865
R348 VSS.t4 VSS.n38 146.865
R349 VSS.t4 VSS.n40 146.865
R350 VSS.t7 VSS.n18 146.865
R351 VSS.t7 VSS.n19 146.865
R352 VSS.n29 VSS.t16 146.865
R353 VSS.n484 VSS.t16 146.865
R354 VSS.n243 VSS.n234 146.505
R355 VSS.n350 VSS.n349 146.25
R356 VSS.n146 VSS.n145 146.25
R357 VSS.n159 VSS.n145 146.25
R358 VSS.n157 VSS.n140 146.25
R359 VSS.n158 VSS.n157 146.25
R360 VSS.n345 VSS.n344 146.25
R361 VSS.n344 VSS.n343 146.25
R362 VSS.n316 VSS.n177 140.8
R363 VSS.n414 VSS.n93 134.489
R364 VSS.n276 VSS.n268 134.489
R365 VSS.n276 VSS.n269 132.659
R366 VSS.n255 VSS.t35 130.689
R367 VSS.n414 VSS.n413 129.781
R368 VSS.n252 VSS.n234 129.781
R369 VSS.n201 VSS.t0 127.005
R370 VSS.n300 VSS.n150 126.721
R371 VSS.n249 VSS.n248 125.746
R372 VSS.n108 VSS.n95 125.365
R373 VSS.n419 VSS.n80 120.484
R374 VSS.n82 VSS.n70 120.484
R375 VSS.n72 VSS.n59 120.484
R376 VSS.n62 VSS.n61 120.484
R377 VSS.n49 VSS.n36 120.484
R378 VSS.n37 VSS.n15 120.484
R379 VSS.n26 VSS.n17 120.484
R380 VSS.n488 VSS.n1 118.416
R381 VSS.n396 VSS.n363 117.379
R382 VSS.n194 VSS.n193 117.001
R383 VSS.n196 VSS.n194 117.001
R384 VSS.n195 VSS.n191 117.001
R385 VSS.n197 VSS.n195 117.001
R386 VSS.n279 VSS.n278 117.001
R387 VSS.n278 VSS.t18 117.001
R388 VSS.n277 VSS.n276 117.001
R389 VSS.t18 VSS.n277 117.001
R390 VSS.n237 VSS.n233 117.001
R391 VSS.n233 VSS.t35 117.001
R392 VSS.n234 VSS.n232 117.001
R393 VSS.n232 VSS.t35 117.001
R394 VSS.n348 VSS.n138 117.001
R395 VSS.n138 VSS.t37 117.001
R396 VSS.n139 VSS.n137 117.001
R397 VSS.n137 VSS.t37 117.001
R398 VSS.n415 VSS.n414 117.001
R399 VSS.n416 VSS.n415 117.001
R400 VSS.n410 VSS.n409 117.001
R401 VSS.n409 VSS.n408 117.001
R402 VSS.n420 VSS.n77 112.942
R403 VSS.n428 VSS.n77 112.942
R404 VSS.n429 VSS.n428 112.942
R405 VSS.n430 VSS.n429 112.942
R406 VSS.n430 VSS.n56 112.942
R407 VSS.n439 VSS.n56 112.942
R408 VSS.n440 VSS.n439 112.942
R409 VSS.n447 VSS.n446 112.942
R410 VSS.n446 VSS.n445 112.942
R411 VSS.n445 VSS.n444 112.942
R412 VSS.n444 VSS.n443 112.942
R413 VSS.n443 VSS.n28 112.942
R414 VSS.n462 VSS.n28 112.942
R415 VSS.n424 VSS.n423 112.942
R416 VSS.n425 VSS.n424 112.942
R417 VSS.n425 VSS.n67 112.942
R418 VSS.n433 VSS.n67 112.942
R419 VSS.n434 VSS.n433 112.942
R420 VSS.n436 VSS.n434 112.942
R421 VSS.n450 VSS.n45 112.942
R422 VSS.n451 VSS.n450 112.942
R423 VSS.n452 VSS.n451 112.942
R424 VSS.n452 VSS.n23 112.942
R425 VSS.n471 VSS.n23 112.942
R426 VSS.n471 VSS.n470 112.942
R427 VSS.n470 VSS.n469 112.942
R428 VSS.n365 VSS.n363 112.93
R429 VSS.n436 VSS.n435 111.436
R430 VSS.n246 VSS.n245 111.112
R431 VSS.n160 VSS.n159 108.213
R432 VSS.n273 VSS.t5 105.689
R433 VSS.n31 VSS.n10 97.4396
R434 VSS.n32 VSS.n12 97.4396
R435 VSS.n372 VSS.n371 97.4396
R436 VSS.n386 VSS.n384 97.4396
R437 VSS.n394 VSS.n393 97.4396
R438 VSS.n377 VSS.n376 96.8664
R439 VSS.n458 VSS.n31 95.7354
R440 VSS.n456 VSS.n32 95.7354
R441 VSS.n371 VSS.n53 95.7354
R442 VSS.n388 VSS.n386 95.7354
R443 VSS.n393 VSS.n390 95.7354
R444 VSS.n376 VSS.n33 95.1723
R445 VSS.n435 VSS.n25 94.352
R446 VSS.n230 VSS.t9 92.5902
R447 VSS.n353 VSS.t9 92.5902
R448 VSS.n406 VSS.n100 91.531
R449 VSS.n461 VSS.n1 87.3879
R450 VSS.n189 VSS.t23 86.7387
R451 VSS.n267 VSS.t19 83.7422
R452 VSS.n121 VSS.t21 83.7278
R453 VSS.n240 VSS.t36 83.7278
R454 VSS.n254 VSS.n231 83.5643
R455 VSS.n404 VSS.n103 82.1622
R456 VSS.n225 VSS.n133 82.1622
R457 VSS.n285 VSS 80.0087
R458 VSS.n245 VSS.t24 77.7783
R459 VSS.n404 VSS.n403 76.5461
R460 VSS.n355 VSS.n133 76.5461
R461 VSS.n114 VSS.n113 76.3709
R462 VSS.n248 VSS.n236 76.3348
R463 VSS.n317 VSS.n176 76.1229
R464 VSS.n305 VSS.n294 75.9791
R465 VSS.n299 VSS.n151 75.6884
R466 VSS.n117 VSS.n108 73.7887
R467 VSS.n204 VSS.n203 73.1255
R468 VSS.n203 VSS.n202 73.1255
R469 VSS.n321 VSS.n169 73.1255
R470 VSS.n169 VSS.n164 73.1255
R471 VSS.n322 VSS.n321 73.1255
R472 VSS.n323 VSS.n322 73.1255
R473 VSS.n175 VSS.n174 73.1255
R474 VSS.n174 VSS.n173 73.1255
R475 VSS.n117 VSS.n116 73.1255
R476 VSS.n116 VSS.n115 73.1255
R477 VSS.n403 VSS.n102 73.1255
R478 VSS.t17 VSS.n102 73.1255
R479 VSS.n103 VSS.n101 73.1255
R480 VSS.t17 VSS.n101 73.1255
R481 VSS.n113 VSS.n95 73.1255
R482 VSS.n285 VSS.n183 73.1255
R483 VSS.n273 VSS.n183 73.1255
R484 VSS.n184 VSS.n182 73.1255
R485 VSS.n294 VSS.n179 73.1255
R486 VSS.n292 VSS.n179 73.1255
R487 VSS.n178 VSS.n177 73.1255
R488 VSS.n291 VSS.n178 73.1255
R489 VSS.n153 VSS.n151 73.1255
R490 VSS.n236 VSS.n228 73.1255
R491 VSS.t24 VSS.n228 73.1255
R492 VSS.n249 VSS.n227 73.1255
R493 VSS.t24 VSS.n227 73.1255
R494 VSS.n355 VSS.n354 73.1255
R495 VSS.n354 VSS.n353 73.1255
R496 VSS.n229 VSS.n225 73.1255
R497 VSS.n230 VSS.n229 73.1255
R498 VSS.n300 VSS.n152 73.1255
R499 VSS.n161 VSS.n152 73.1255
R500 VSS.n147 VSS.n146 71.5299
R501 VSS.n289 VSS.n288 65.232
R502 VSS.n408 VSS.n407 64.8941
R503 VSS.n351 VSS.t25 63.4558
R504 VSS.n329 VSS.n161 62.5456
R505 VSS.n220 VSS.n184 62.3981
R506 VSS.n486 VSS.n485 62.305
R507 VSS.n465 VSS.n25 61.8241
R508 VSS.n447 VSS.n441 61.7417
R509 VSS.n482 VSS.n481 61.2169
R510 VSS.n407 VSS.n406 59.6587
R511 VSS.t38 VSS.n418 58.6566
R512 VSS.t38 VSS.n419 58.6566
R513 VSS.t8 VSS.n80 58.6566
R514 VSS.t8 VSS.n82 58.6566
R515 VSS.t6 VSS.n70 58.6566
R516 VSS.t6 VSS.n72 58.6566
R517 VSS.t10 VSS.n59 58.6566
R518 VSS.t10 VSS.n62 58.6566
R519 VSS.t11 VSS.n49 58.6566
R520 VSS.t4 VSS.n36 58.6566
R521 VSS.t4 VSS.n37 58.6566
R522 VSS.t7 VSS.n15 58.6566
R523 VSS.t7 VSS.n17 58.6566
R524 VSS.n26 VSS.t16 58.6566
R525 VSS.n466 VSS.t16 58.6566
R526 VSS.t32 VSS.n5 58.6566
R527 VSS.t24 VSS.t35 58.2016
R528 VSS.n408 VSS.t20 56.0289
R529 VSS.n416 VSS.t20 56.0289
R530 VSS.n293 VSS.n292 55.0005
R531 VSS.n206 VSS.n192 54.9719
R532 VSS.n150 VSS.n147 53.3135
R533 VSS.n441 VSS.n440 51.2005
R534 VSS.n462 VSS.n461 49.3181
R535 VSS.n469 VSS.n25 49.3181
R536 VSS.n369 VSS.n50 48.6248
R537 VSS.n482 VSS.n9 47.5841
R538 VSS.n333 VSS.n332 46.3872
R539 VSS.n280 VSS.n268 43.5902
R540 VSS.n199 VSS.n198 41.7862
R541 VSS.t0 VSS.n199 41.7862
R542 VSS.n172 VSS.n166 41.7862
R543 VSS.t28 VSS.n166 41.7862
R544 VSS.n200 VSS.n170 41.7862
R545 VSS.t0 VSS.n200 41.7862
R546 VSS.n319 VSS.n167 41.7862
R547 VSS.t28 VSS.n167 41.7862
R548 VSS.n309 VSS.n308 41.7862
R549 VSS.n308 VSS.t2 41.7862
R550 VSS.n307 VSS.n306 41.7862
R551 VSS.t2 VSS.n307 41.7862
R552 VSS.n334 VSS.n333 41.7862
R553 VSS.n304 VSS.n303 41.7862
R554 VSS.n303 VSS.n302 41.7862
R555 VSS.n188 VSS.t1 41.7156
R556 VSS.n295 VSS.t3 41.4575
R557 VSS.n297 VSS.t31 41.4563
R558 VSS.n311 VSS.t29 41.4498
R559 VSS.n279 VSS.n269 39.8737
R560 VSS.n213 VSS.n190 39.1319
R561 VSS.n213 VSS.n191 38.7101
R562 VSS.n246 VSS.n154 38.6075
R563 VSS.n210 VSS.n193 37.7441
R564 VSS.n352 VSS.n351 37.2102
R565 VSS.n115 VSS.n112 36.7801
R566 VSS.n290 VSS.n165 36.2505
R567 VSS.n298 VSS.n149 34.0553
R568 VSS.n210 VSS.n209 32.9148
R569 VSS.n242 VSS.n241 32.377
R570 VSS.n242 VSS.n235 30.1719
R571 VSS.n353 VSS.n352 30.1064
R572 VSS.t11 VSS.n50 28.0386
R573 VSS.n305 VSS.n299 26.3819
R574 VSS.n417 VSS.n416 25.1778
R575 VSS.n342 VSS.n341 23.4005
R576 VSS.n342 VSS.t25 23.4005
R577 VSS.n144 VSS.n142 23.4005
R578 VSS.n144 VSS.t25 23.4005
R579 VSS.n176 VSS.n175 21.7605
R580 VSS.n211 VSS.n192 19.81
R581 VSS.n61 VSS.n50 19.4204
R582 VSS.n264 VSS.n222 18.5973
R583 VSS.n403 VSS 17.8552
R584 VSS VSS.n355 17.8552
R585 VSS.n220 VSS.n185 17.4457
R586 VSS.n481 VSS.n480 16.8875
R587 VSS.n309 VSS.n149 16.6656
R588 VSS.n413 VSS.n412 16.5348
R589 VSS.n206 VSS.n205 16.4078
R590 VSS.n96 VSS.n93 16.4078
R591 VSS.n335 VSS.n149 16.3973
R592 VSS.n460 VSS.n9 16.2503
R593 VSS.n481 VSS.n479 15.2441
R594 VSS.n474 VSS.n12 15.2441
R595 VSS.n373 VSS.n12 15.2441
R596 VSS.n378 VSS.n377 15.2441
R597 VSS.n372 VSS.n367 15.2441
R598 VSS.n384 VSS.n383 15.2441
R599 VSS.n395 VSS.n394 15.2441
R600 VSS.n478 VSS.n10 14.7787
R601 VSS.n384 VSS.n382 14.7787
R602 VSS.n394 VSS.n364 14.7787
R603 VSS.n475 VSS.n10 14.546
R604 VSS.n377 VSS.n374 14.546
R605 VSS.n112 VSS.n99 14.5188
R606 VSS.n118 VSS.n107 14.2116
R607 VSS.n379 VSS.n372 13.615
R608 VSS.n118 VSS.n117 13.4459
R609 VSS.n243 VSS.n242 13.1205
R610 VSS.n54 VSS.n33 12.4289
R611 VSS.n390 VSS.n365 12.3876
R612 VSS.n390 VSS.n389 12.3876
R613 VSS.n389 VSS.n388 12.3876
R614 VSS.n388 VSS.n387 12.3876
R615 VSS.n387 VSS.n53 12.3876
R616 VSS.n456 VSS.n455 12.3876
R617 VSS.n457 VSS.n456 12.3876
R618 VSS.n458 VSS.n457 12.3876
R619 VSS.n459 VSS.n458 12.3876
R620 VSS.n455 VSS.n33 12.3463
R621 VSS.n411 VSS.n96 11.8862
R622 VSS.n465 VSS.n464 11.6307
R623 VSS.n128 VSS.n106 11.6134
R624 VSS.n260 VSS.n224 11.6134
R625 VSS.n321 VSS.n168 11.5469
R626 VSS.n321 VSS.n320 11.217
R627 VSS.n236 VSS.n222 10.7568
R628 VSS.n252 VSS.n251 10.4904
R629 VSS.n315 VSS.n310 10.4191
R630 VSS.n345 VSS.n143 10.2128
R631 VSS.n292 VSS.n154 10.0005
R632 VSS.n193 VSS.n192 9.84665
R633 VSS.n120 VSS.n118 9.41534
R634 VSS.n261 VSS.n260 9.39185
R635 VSS.n212 VSS.n211 9.37653
R636 VSS.n346 VSS.n345 9.3005
R637 VSS.n221 VSS.n220 9.3005
R638 VSS.n129 VSS.n128 9.3005
R639 VSS.n412 VSS.n94 9.06717
R640 VSS.n386 VSS.n366 8.0142
R641 VSS.n366 VSS.n75 8.0142
R642 VSS.n371 VSS.n368 8.0142
R643 VSS.n368 VSS.n65 8.0142
R644 VSS.n386 VSS.n385 8.0142
R645 VSS.n385 VSS.n63 8.0142
R646 VSS.n376 VSS.n375 8.0142
R647 VSS.n375 VSS.n52 8.0142
R648 VSS.n371 VSS.n370 8.0142
R649 VSS.n370 VSS.n369 8.0142
R650 VSS.n35 VSS.n32 8.0142
R651 VSS.n40 VSS.n35 8.0142
R652 VSS.n376 VSS.n34 8.0142
R653 VSS.n38 VSS.n34 8.0142
R654 VSS.n31 VSS.n14 8.0142
R655 VSS.n19 VSS.n14 8.0142
R656 VSS.n32 VSS.n13 8.0142
R657 VSS.n18 VSS.n13 8.0142
R658 VSS.n31 VSS.n30 8.0142
R659 VSS.n30 VSS.n29 8.0142
R660 VSS.n393 VSS.n391 8.0142
R661 VSS.n391 VSS.n85 8.0142
R662 VSS.n393 VSS.n392 8.0142
R663 VSS.n392 VSS.n73 8.0142
R664 VSS.n363 VSS.n362 8.0142
R665 VSS.n362 VSS.n83 8.0142
R666 VSS.n483 VSS.n482 8.0142
R667 VSS.n484 VSS.n483 8.0142
R668 VSS.n340 VSS.n143 7.99658
R669 VSS.n412 VSS.n95 7.60521
R670 VSS.t5 VSS.n181 7.50192
R671 VSS.n128 VSS.n127 7.48437
R672 VSS.n260 VSS.n259 7.48437
R673 VSS.n341 VSS.n147 7.45136
R674 VSS.n489 VSS.n0 7.30675
R675 VSS.n211 VSS.n210 7.13193
R676 VSS.n106 VSS.n104 6.92198
R677 VSS.n224 VSS.n132 6.92198
R678 VSS.n441 VSS.n54 6.77211
R679 VSS.n347 VSS.n346 6.74718
R680 VSS.n205 VSS.n204 6.4257
R681 VSS.n412 VSS.n411 6.4005
R682 VSS.n320 VSS.n170 6.18574
R683 VSS.n320 VSS.n319 6.18574
R684 VSS VSS.n489 5.91834
R685 VSS.n441 VSS.n53 5.61598
R686 VSS VSS.n284 5.45235
R687 VSS VSS.n402 5.45235
R688 VSS.n356 VSS 5.45235
R689 VSS.n127 VSS.n103 5.41985
R690 VSS.n259 VSS.n225 5.41985
R691 VSS.n460 VSS.n459 5.40953
R692 VSS.n255 VSS.n254 5.29151
R693 VSS.n161 VSS.n160 4.9644
R694 VSS VSS.n222 4.92986
R695 VSS.n214 VSS.n213 4.90573
R696 VSS.n318 VSS.n317 4.59111
R697 VSS.n89 VSS.n86 4.46615
R698 VSS.n419 VSS.n89 4.46615
R699 VSS.n79 VSS.n76 4.46615
R700 VSS.n82 VSS.n79 4.46615
R701 VSS.n86 VSS.n78 4.46615
R702 VSS.n80 VSS.n78 4.46615
R703 VSS.n69 VSS.n66 4.46615
R704 VSS.n72 VSS.n69 4.46615
R705 VSS.n76 VSS.n68 4.46615
R706 VSS.n70 VSS.n68 4.46615
R707 VSS.n58 VSS.n55 4.46615
R708 VSS.n62 VSS.n58 4.46615
R709 VSS.n66 VSS.n57 4.46615
R710 VSS.n59 VSS.n57 4.46615
R711 VSS.n47 VSS.n44 4.46615
R712 VSS.n49 VSS.n47 4.46615
R713 VSS.n55 VSS.n46 4.46615
R714 VSS.n61 VSS.n46 4.46615
R715 VSS.n442 VSS.n43 4.46615
R716 VSS.n43 VSS.n37 4.46615
R717 VSS.n44 VSS.n42 4.46615
R718 VSS.n42 VSS.n36 4.46615
R719 VSS.n24 VSS.n22 4.46615
R720 VSS.n22 VSS.n17 4.46615
R721 VSS.n442 VSS.n21 4.46615
R722 VSS.n21 VSS.n15 4.46615
R723 VSS.n27 VSS.n24 4.46615
R724 VSS.n27 VSS.n26 4.46615
R725 VSS.n88 VSS.n87 4.46615
R726 VSS.n418 VSS.n88 4.46615
R727 VSS.n467 VSS.n465 4.46615
R728 VSS.n467 VSS.n466 4.46615
R729 VSS.n9 VSS.n8 4.46615
R730 VSS.n8 VSS.n5 4.46615
R731 VSS.n487 VSS.n486 4.46615
R732 VSS.n251 VSS.n250 4.44728
R733 VSS.n298 VSS.n294 4.36414
R734 VSS.n259 VSS.n226 4.35795
R735 VSS.n461 VSS.n460 4.09269
R736 VSS.n398 VSS.n397 3.87676
R737 VSS.n250 VSS.n249 3.8405
R738 VSS VSS.n94 3.37828
R739 VSS.n215 VSS.n170 3.29929
R740 VSS.t17 VSS.n114 3.10271
R741 VSS.n298 VSS.n295 3.1005
R742 VSS.n298 VSS.n297 3.1005
R743 VSS.n250 VSS.n226 2.86007
R744 VSS.n284 VSS.n283 2.3255
R745 VSS.n125 VSS.n124 2.3255
R746 VSS.n402 VSS.n401 2.3255
R747 VSS.n357 VSS.n356 2.3255
R748 VSS.n258 VSS.n223 2.3255
R749 VSS.n126 VSS 2.31161
R750 VSS.n257 VSS 2.28816
R751 VSS.n251 VSS.n235 2.13383
R752 VSS.n190 VSS.n189 1.89317
R753 VSS.n121 VSS.n97 1.86348
R754 VSS.n241 VSS.n240 1.86348
R755 VSS.n311 VSS.n176 1.8605
R756 VSS.n214 VSS.n188 1.8605
R757 VSS.n364 VSS.n361 1.8605
R758 VSS.n382 VSS.n381 1.8605
R759 VSS.n380 VSS.n379 1.8605
R760 VSS.n374 VSS.n11 1.8605
R761 VSS.n476 VSS.n475 1.8605
R762 VSS.n478 VSS.n477 1.8605
R763 VSS.n281 VSS.n280 1.8605
R764 VSS.n397 VSS.n396 1.8605
R765 VSS.n317 VSS.n316 1.85321
R766 VSS.n126 VSS.n125 1.77828
R767 VSS.n213 VSS.n212 1.66708
R768 VSS.n398 VSS.n360 1.64434
R769 VSS.n379 VSS.n378 1.62959
R770 VSS.n127 VSS.n126 1.61889
R771 VSS.n435 VSS.n45 1.50638
R772 VSS.n299 VSS.n298 1.46981
R773 VSS.n259 VSS.n258 1.3622
R774 VSS.n123 VSS.n94 1.32907
R775 VSS.n238 VSS.n226 1.32907
R776 VSS.n348 VSS.n347 1.2805
R777 VSS.n337 VSS 1.2505
R778 VSS.n359 VSS 1.2505
R779 VSS.n186 VSS.t12 1.21428
R780 VSS.t15 VSS.n219 1.21428
R781 VSS.n411 VSS.n410 1.20521
R782 VSS.n237 VSS.n235 1.20521
R783 VSS.n312 VSS.n311 1.06892
R784 VSS.n219 VSS.n186 1.04896
R785 VSS.n204 VSS.n191 1.00837
R786 VSS VSS.n265 0.976194
R787 VSS.n400 VSS.n129 0.971333
R788 VSS.n221 VSS.t15 0.909702
R789 VSS.n477 VSS 0.896681
R790 VSS.n313 VSS.n310 0.845955
R791 VSS.n336 VSS.n335 0.845955
R792 VSS.n475 VSS.n474 0.698682
R793 VSS.n485 VSS.t32 0.673635
R794 VSS.n318 VSS.n171 0.592183
R795 VSS.n340 VSS.n339 0.529939
R796 VSS.n217 VSS.n171 0.520386
R797 VSS.n216 VSS.n215 0.517167
R798 VSS.n143 VSS.n141 0.517167
R799 VSS.n212 VSS.n187 0.517167
R800 VSS.t14 VSS.n218 0.473714
R801 VSS.n479 VSS.n478 0.465955
R802 VSS.n374 VSS.n373 0.465955
R803 VSS.n382 VSS.n367 0.465955
R804 VSS.n383 VSS.n364 0.465955
R805 VSS.n396 VSS.n395 0.465955
R806 VSS.n339 VSS.n336 0.462148
R807 VSS.n280 VSS.n279 0.457643
R808 VSS.n2 VSS.n0 0.436436
R809 VSS.n358 VSS.n130 0.407111
R810 VSS.n346 VSS.n141 0.405672
R811 VSS.n97 VSS.n96 0.376971
R812 VSS.n283 VSS.n282 0.367087
R813 VSS.n399 VSS.n398 0.360165
R814 VSS.n119 VSS.n106 0.321176
R815 VSS.n123 VSS.n122 0.320051
R816 VSS.n262 VSS.n224 0.315718
R817 VSS.n360 VSS.n358 0.296949
R818 VSS.n310 VSS.n309 0.268407
R819 VSS.n335 VSS.n334 0.268407
R820 VSS.n239 VSS.n238 0.263801
R821 VSS.n490 VSS 0.2605
R822 VSS.n339 VSS 0.236295
R823 VSS VSS.n357 0.232471
R824 VSS.n464 VSS.n1 0.231743
R825 VSS.n218 VSS.n217 0.21925
R826 VSS.n399 VSS 0.216846
R827 VSS.n380 VSS.n11 0.212306
R828 VSS.n476 VSS.n11 0.212306
R829 VSS.n397 VSS.n361 0.208833
R830 VSS.n381 VSS.n361 0.208833
R831 VSS.n381 VSS.n380 0.205361
R832 VSS.n477 VSS.n476 0.205361
R833 VSS.n240 VSS.n239 0.197673
R834 VSS.n338 VSS.n141 0.194466
R835 VSS.n341 VSS.n340 0.188758
R836 VSS.n209 VSS.n190 0.183357
R837 VSS.n490 VSS.n0 0.18175
R838 VSS.n263 VSS.n223 0.176839
R839 VSS.n265 VSS.n264 0.172797
R840 VSS.n313 VSS.n148 0.172375
R841 VSS.n336 VSS.n148 0.166693
R842 VSS.n186 VSS.t13 0.165823
R843 VSS.n219 VSS.t14 0.165823
R844 VSS.n216 VSS.n188 0.163852
R845 VSS.n131 VSS.n130 0.152527
R846 VSS.n189 VSS.n187 0.151068
R847 VSS.n296 VSS.n148 0.146333
R848 VSS.n120 VSS.n119 0.143095
R849 VSS.n312 VSS.n171 0.141125
R850 VSS.n218 VSS.n187 0.136864
R851 VSS.n217 VSS.n216 0.128341
R852 VSS.n401 VSS.n105 0.1255
R853 VSS.n314 VSS.n312 0.122659
R854 VSS.n122 VSS.n121 0.119548
R855 VSS.n266 VSS 0.113
R856 VSS.n263 VSS.n262 0.10958
R857 VSS.n265 VSS.n130 0.108139
R858 VSS.n490 VSS 0.105518
R859 VSS.n338 VSS.n337 0.0999318
R860 VSS.n314 VSS.n313 0.0999318
R861 VSS.n124 VSS.n123 0.0954519
R862 VSS.n238 VSS.n223 0.0954519
R863 VSS.n267 VSS.n266 0.0934487
R864 VSS VSS.n281 0.088641
R865 VSS.n264 VSS.n263 0.0861481
R866 VSS.n358 VSS 0.0835761
R867 VSS.n129 VSS.n105 0.0796667
R868 VSS.n319 VSS.n318 0.0729516
R869 VSS.n360 VSS.n359 0.0714459
R870 VSS.n122 VSS 0.06925
R871 VSS.n283 VSS.n221 0.0684987
R872 VSS.n357 VSS.n131 0.063
R873 VSS.n124 VSS.n120 0.0593663
R874 VSS VSS.n338 0.0558977
R875 VSS VSS.n490 0.05425
R876 VSS.n261 VSS.n131 0.0540714
R877 VSS.n410 VSS.n97 0.0506961
R878 VSS.n241 VSS.n237 0.0506961
R879 VSS.n489 VSS.n488 0.0481923
R880 VSS.n284 VSS.n185 0.0479074
R881 VSS.n402 VSS.n104 0.0479074
R882 VSS.n356 VSS.n132 0.0479074
R883 VSS.n239 VSS 0.047375
R884 VSS.n315 VSS.n314 0.047
R885 VSS.n215 VSS.n214 0.043453
R886 VSS.n282 VSS 0.0402727
R887 VSS.n125 VSS.n107 0.0360556
R888 VSS.n266 VSS 0.0325513
R889 VSS.n296 VSS.n295 0.03175
R890 VSS.n297 VSS.n296 0.03175
R891 VSS.n258 VSS.n257 0.027734
R892 VSS.n282 VSS 0.0229359
R893 VSS.n262 VSS.n261 0.0192927
R894 VSS.n119 VSS.n105 0.0180921
R895 VSS.n401 VSS.n400 0.0125192
R896 VSS.n400 VSS.n399 0.0101154
R897 VSS.n359 VSS 0.00387838
R898 VSS.n337 VSS 0.00334091
R899 VSS.n281 VSS.n267 0.00210256
R900 x1.x1.pg2g x1.x1.pg2g.t1 61.169
R901 x1.x1.pg2g x1.x1.pg2g.t2 22.3222
R902 x1.x1.pg2g x1.x1.pg2g.t0 21.7234
R903 x1.x1.mirhigh.n0 x1.x1.mirhigh.t0 73.9922
R904 x1.x1.mirhigh x1.x1.mirhigh.t1 62.3033
R905 x1.x1.mirhigh.n0 x1.x1.mirhigh.t2 48.1635
R906 x1.x1.mirhigh x1.x1.mirhigh.n0 1.99219
R907 VCC.n88 VCC.n87 4560
R908 VCC.n85 VCC.n83 4560
R909 VCC.n73 VCC.n70 4560
R910 VCC.n76 VCC.n69 4560
R911 VCC.n34 VCC.n32 4560
R912 VCC.n37 VCC.n36 4560
R913 VCC.n102 VCC.n15 4207.06
R914 VCC.n99 VCC.n16 4207.06
R915 VCC.n49 VCC.n43 3854.12
R916 VCC.n47 VCC.n46 3854.12
R917 VCC.n26 VCC.n25 3854.12
R918 VCC.n23 VCC.n21 3854.12
R919 VCC.n62 VCC.n56 2848.24
R920 VCC.n60 VCC.n59 2848.24
R921 VCC.n216 VCC.n210 1860
R922 VCC.n213 VCC.n211 1860
R923 VCC.n161 VCC.n155 1860
R924 VCC.n159 VCC.n158 1860
R925 VCC.n145 VCC.n139 1860
R926 VCC.n143 VCC.n142 1860
R927 VCC.n189 VCC.n183 1807.06
R928 VCC.n186 VCC.n184 1807.06
R929 VCC.n199 VCC.n197 1807.06
R930 VCC.n202 VCC.n196 1807.06
R931 VCC.n130 VCC.n123 1807.06
R932 VCC.n127 VCC.n124 1807.06
R933 VCC.n115 VCC.n108 1807.06
R934 VCC.n112 VCC.n109 1807.06
R935 VCC.n176 VCC.n169 1807.06
R936 VCC.n173 VCC.n170 1807.06
R937 VCC.n9 VCC.n8 1736.47
R938 VCC.n6 VCC.n4 1736.47
R939 VCC.n100 VCC.n15 1068.61
R940 VCC.n101 VCC.n16 1068.61
R941 VCC.n59 VCC.n58 1018.62
R942 VCC.n62 VCC.n61 1018.62
R943 VCC.n74 VCC.n69 879.971
R944 VCC.n75 VCC.n70 879.971
R945 VCC.n200 VCC.n196 594.523
R946 VCC.n201 VCC.n197 594.523
R947 VCC.n113 VCC.n112 594.523
R948 VCC.n115 VCC.n114 594.523
R949 VCC.n158 VCC.n157 561.481
R950 VCC.n161 VCC.n160 561.481
R951 VCC.n142 VCC.n141 561.481
R952 VCC.n145 VCC.n144 561.481
R953 VCC.n84 VCC.n80 486.401
R954 VCC.n84 VCC.n81 486.401
R955 VCC.n89 VCC.n81 486.401
R956 VCC.n77 VCC.n68 486.401
R957 VCC.n33 VCC.n29 486.401
R958 VCC.n33 VCC.n30 486.401
R959 VCC.n38 VCC.n30 486.401
R960 VCC.n78 VCC.n77 468.406
R961 VCC.n103 VCC.n14 443.728
R962 VCC.n104 VCC.n103 436.236
R963 VCC.n50 VCC.n42 411.106
R964 VCC.n44 VCC.n42 411.106
R965 VCC.n22 VCC.n18 411.106
R966 VCC.n22 VCC.n19 411.106
R967 VCC.n44 VCC.n41 387.128
R968 VCC.n46 VCC.n45 385.567
R969 VCC.n49 VCC.n48 385.567
R970 VCC.n26 VCC.n20 385.567
R971 VCC.n24 VCC.n23 385.567
R972 VCC.n51 VCC.n50 384.087
R973 VCC.n27 VCC.n19 354.171
R974 VCC.n72 VCC.n67 349.312
R975 VCC.n71 VCC.n68 333.82
R976 VCC.n28 VCC.n18 321.255
R977 VCC.n9 VCC.n3 314.781
R978 VCC.n7 VCC.n6 314.781
R979 VCC.n63 VCC.n55 303.812
R980 VCC.n57 VCC.n55 303.812
R981 VCC.n98 VCC.n17 285.354
R982 VCC.n97 VCC.n13 272.99
R983 VCC.n90 VCC.n89 265.865
R984 VCC.n39 VCC.n29 249.901
R985 VCC.n91 VCC.t12 228.284
R986 VCC.n57 VCC.n54 215.555
R987 VCC.n64 VCC.n63 213.397
R988 VCC.n212 VCC.n209 198.4
R989 VCC.n217 VCC.n209 198.4
R990 VCC.n162 VCC.n154 198.4
R991 VCC.n156 VCC.n154 198.4
R992 VCC.n146 VCC.n138 198.4
R993 VCC.n140 VCC.n138 198.4
R994 VCC.n214 VCC.n210 194.888
R995 VCC.n215 VCC.n211 194.888
R996 VCC.n190 VCC.n182 192.754
R997 VCC.n185 VCC.n182 192.754
R998 VCC.n203 VCC.n195 192.754
R999 VCC.n198 VCC.n195 192.754
R1000 VCC.n131 VCC.n122 192.754
R1001 VCC.n126 VCC.n122 192.754
R1002 VCC.n111 VCC.n110 192.754
R1003 VCC.n111 VCC.n106 192.754
R1004 VCC.n177 VCC.n168 192.754
R1005 VCC.n172 VCC.n168 192.754
R1006 VCC.n90 VCC.n80 186.805
R1007 VCC.n39 VCC.n38 185.901
R1008 VCC.n5 VCC.n1 185.225
R1009 VCC.n5 VCC.n2 185.225
R1010 VCC.n189 VCC.n188 178.274
R1011 VCC.n187 VCC.n186 178.274
R1012 VCC.n130 VCC.n129 178.274
R1013 VCC.n128 VCC.n127 178.274
R1014 VCC.n176 VCC.n175 178.274
R1015 VCC.n174 VCC.n173 178.274
R1016 VCC.n212 VCC.n208 175.391
R1017 VCC.n156 VCC.n153 175.391
R1018 VCC.n140 VCC.n137 175.391
R1019 VCC.n218 VCC.n217 173.403
R1020 VCC.n163 VCC.n162 173.403
R1021 VCC.n147 VCC.n146 173.403
R1022 VCC.n10 VCC.n2 162.456
R1023 VCC.n88 VCC.n82 160.32
R1024 VCC.n86 VCC.n85 160.32
R1025 VCC.n35 VCC.n34 160.32
R1026 VCC.n37 VCC.n31 160.32
R1027 VCC.n11 VCC.n1 159.474
R1028 VCC.n191 VCC.n190 141.655
R1029 VCC.n204 VCC.n203 141.655
R1030 VCC.n132 VCC.n131 141.655
R1031 VCC.n117 VCC.n106 141.655
R1032 VCC.n178 VCC.n177 141.655
R1033 VCC.n79 VCC.t3 113.716
R1034 VCC.n136 VCC.t8 113.68
R1035 VCC.n220 VCC.t10 113.644
R1036 VCC.n152 VCC.t1 113.644
R1037 VCC.n183 VCC.n181 92.5005
R1038 VCC.n184 VCC.n182 92.5005
R1039 VCC.n197 VCC.n194 92.5005
R1040 VCC.n196 VCC.n195 92.5005
R1041 VCC.n123 VCC.n121 92.5005
R1042 VCC.n124 VCC.n122 92.5005
R1043 VCC.n112 VCC.n111 92.5005
R1044 VCC.n116 VCC.n115 92.5005
R1045 VCC.n169 VCC.n167 92.5005
R1046 VCC.n170 VCC.n168 92.5005
R1047 VCC.n63 VCC.n62 92.5005
R1048 VCC.n59 VCC.n57 92.5005
R1049 VCC.n187 VCC.n183 79.3155
R1050 VCC.n188 VCC.n184 79.3155
R1051 VCC.n128 VCC.n123 79.3155
R1052 VCC.n129 VCC.n124 79.3155
R1053 VCC.n174 VCC.n169 79.3155
R1054 VCC.n175 VCC.n170 79.3155
R1055 VCC.n185 VCC.n180 72.9076
R1056 VCC.n198 VCC.n193 72.9076
R1057 VCC.n126 VCC.n125 72.9076
R1058 VCC.n110 VCC.n107 72.9076
R1059 VCC.n172 VCC.n171 72.9076
R1060 VCC.n213 VCC.n212 61.6672
R1061 VCC.n217 VCC.n216 61.6672
R1062 VCC.n162 VCC.n161 61.6672
R1063 VCC.n158 VCC.n156 61.6672
R1064 VCC.n146 VCC.n145 61.6672
R1065 VCC.n142 VCC.n140 61.6672
R1066 VCC.n214 VCC.n213 53.4348
R1067 VCC.n216 VCC.n215 53.4348
R1068 VCC.n53 VCC.t19 48.1635
R1069 VCC.n4 VCC.n1 37.0005
R1070 VCC.n8 VCC.n2 37.0005
R1071 VCC.n16 VCC.n14 30.8338
R1072 VCC.n15 VCC.n13 30.8338
R1073 VCC.n6 VCC.n5 30.8338
R1074 VCC.n10 VCC.n9 30.8338
R1075 VCC.n4 VCC.n3 29.6618
R1076 VCC.n8 VCC.n7 29.6618
R1077 VCC.n190 VCC.n189 23.1255
R1078 VCC.n186 VCC.n185 23.1255
R1079 VCC.n211 VCC.n209 23.1255
R1080 VCC.n210 VCC.n208 23.1255
R1081 VCC.n203 VCC.n202 23.1255
R1082 VCC.n199 VCC.n198 23.1255
R1083 VCC.n159 VCC.n154 23.1255
R1084 VCC.n155 VCC.n153 23.1255
R1085 VCC.n131 VCC.n130 23.1255
R1086 VCC.n127 VCC.n126 23.1255
R1087 VCC.n143 VCC.n138 23.1255
R1088 VCC.n139 VCC.n137 23.1255
R1089 VCC.n110 VCC.n109 23.1255
R1090 VCC.n108 VCC.n106 23.1255
R1091 VCC.n177 VCC.n176 23.1255
R1092 VCC.n173 VCC.n172 23.1255
R1093 VCC.n83 VCC.n80 23.1255
R1094 VCC.n87 VCC.n81 23.1255
R1095 VCC.n70 VCC.n67 23.1255
R1096 VCC.n69 VCC.n68 23.1255
R1097 VCC.n32 VCC.n29 23.1255
R1098 VCC.n36 VCC.n30 23.1255
R1099 VCC.n83 VCC.n82 22.2004
R1100 VCC.n87 VCC.n86 22.2004
R1101 VCC.n32 VCC.n31 22.2004
R1102 VCC.n36 VCC.n35 22.2004
R1103 VCC.n181 VCC.n180 21.8808
R1104 VCC.n194 VCC.n193 21.8808
R1105 VCC.n125 VCC.n121 21.8808
R1106 VCC.n116 VCC.n107 21.8808
R1107 VCC.n171 VCC.n167 21.8808
R1108 VCC.n157 VCC.n155 15.947
R1109 VCC.n160 VCC.n159 15.947
R1110 VCC.n141 VCC.n139 15.947
R1111 VCC.n144 VCC.n143 15.947
R1112 VCC.n200 VCC.n199 15.3218
R1113 VCC.n202 VCC.n201 15.3218
R1114 VCC.n113 VCC.n108 15.3218
R1115 VCC.n114 VCC.n109 15.3218
R1116 VCC.n50 VCC.n49 13.2148
R1117 VCC.n47 VCC.n42 13.2148
R1118 VCC.n46 VCC.n44 13.2148
R1119 VCC.n43 VCC.n41 13.2148
R1120 VCC.n21 VCC.n18 13.2148
R1121 VCC.n23 VCC.n22 13.2148
R1122 VCC.n25 VCC.n19 13.2148
R1123 VCC.n27 VCC.n26 13.2148
R1124 VCC.n28 VCC.n27 13.0138
R1125 VCC.n45 VCC.n43 11.8527
R1126 VCC.n48 VCC.n47 11.8527
R1127 VCC.n21 VCC.n20 11.8527
R1128 VCC.n25 VCC.n24 11.8527
R1129 VCC.n60 VCC.n55 10.8829
R1130 VCC.n56 VCC.n54 10.8829
R1131 VCC.n125 VCC.n120 10.0831
R1132 VCC.n192 VCC.n180 9.48305
R1133 VCC.n107 VCC 9.44764
R1134 VCC.n206 VCC.n193 9.37472
R1135 VCC.n171 VCC.n166 9.37472
R1136 VCC.t4 VCC.n187 9.12649
R1137 VCC.n188 VCC.t4 9.12649
R1138 VCC.t5 VCC.n128 9.12649
R1139 VCC.n129 VCC.t5 9.12649
R1140 VCC.t20 VCC.n174 9.12649
R1141 VCC.n175 VCC.t20 9.12649
R1142 VCC.n72 VCC.n71 9.08437
R1143 VCC.n12 VCC.t22 8.96809
R1144 VCC.n201 VCC.t6 7.60912
R1145 VCC.t6 VCC.n200 7.60912
R1146 VCC.n114 VCC.t14 7.60912
R1147 VCC.t14 VCC.n113 7.60912
R1148 VCC.n77 VCC.n76 7.4005
R1149 VCC.n73 VCC.n72 7.4005
R1150 VCC.n99 VCC.n98 7.4005
R1151 VCC.n103 VCC.n102 7.4005
R1152 VCC.n85 VCC.n84 7.11588
R1153 VCC.n89 VCC.n88 7.11588
R1154 VCC.n34 VCC.n33 7.11588
R1155 VCC.n38 VCC.n37 7.11588
R1156 VCC VCC.n95 7.00201
R1157 VCC.n160 VCC.t0 6.98177
R1158 VCC.n157 VCC.t0 6.98177
R1159 VCC.n144 VCC.t7 6.98177
R1160 VCC.n141 VCC.t7 6.98177
R1161 VCC.n58 VCC.n56 6.96486
R1162 VCC.n61 VCC.n60 6.96486
R1163 VCC.n7 VCC.t13 6.70818
R1164 VCC.t13 VCC.n3 6.70818
R1165 VCC.n215 VCC.t9 6.46232
R1166 VCC.t9 VCC.n214 6.46232
R1167 VCC.n74 VCC.n73 5.9633
R1168 VCC.n76 VCC.n75 5.9633
R1169 VCC.n100 VCC.n99 5.51167
R1170 VCC.n102 VCC.n101 5.51167
R1171 VCC.n78 VCC.n67 4.8645
R1172 VCC.n61 VCC.t18 3.89288
R1173 VCC.n58 VCC.t18 3.89288
R1174 VCC.n52 VCC.n40 3.72362
R1175 VCC.n79 VCC.n78 3.1005
R1176 VCC.n91 VCC.n17 3.1005
R1177 VCC.n95 VCC 2.8755
R1178 VCC.n98 VCC.n97 2.84494
R1179 VCC.n92 VCC.n90 2.6261
R1180 VCC.n222 VCC.n221 2.60004
R1181 VCC.n192 VCC.n191 2.3255
R1182 VCC.n205 VCC.n204 2.3255
R1183 VCC.n133 VCC.n132 2.3255
R1184 VCC.n118 VCC.n117 2.3255
R1185 VCC.n179 VCC.n178 2.3255
R1186 VCC.n52 VCC.n51 1.9301
R1187 VCC.n17 VCC.n14 1.9205
R1188 VCC.n101 VCC.t11 1.88064
R1189 VCC.t11 VCC.n100 1.88064
R1190 VCC.n219 VCC.n218 1.8605
R1191 VCC.n148 VCC.n147 1.8605
R1192 VCC.n164 VCC.n163 1.8605
R1193 VCC.n12 VCC.n11 1.8605
R1194 VCC.n105 VCC.n104 1.8605
R1195 VCC.n40 VCC.n39 1.663
R1196 VCC.n223 VCC.n222 1.56691
R1197 VCC.n11 VCC.n10 1.5365
R1198 VCC.n51 VCC.n41 1.47742
R1199 VCC.n75 VCC.t2 1.42902
R1200 VCC.t2 VCC.n74 1.42902
R1201 VCC.n48 VCC.t16 1.32296
R1202 VCC.n45 VCC.t16 1.32296
R1203 VCC.n24 VCC.t17 1.32296
R1204 VCC.t17 VCC.n20 1.32296
R1205 VCC.n221 VCC.n220 1.31592
R1206 VCC.n104 VCC.n13 1.2805
R1207 VCC.n151 VCC.n118 1.08528
R1208 VCC.n218 VCC.n208 1.0245
R1209 VCC.n163 VCC.n153 1.0245
R1210 VCC.n147 VCC.n137 1.0245
R1211 VCC.n152 VCC.n151 0.915511
R1212 VCC.n64 VCC.n54 0.853833
R1213 VCC.n40 VCC.n28 0.846486
R1214 VCC.n221 VCC 0.839158
R1215 VCC.n86 VCC.t21 0.814017
R1216 VCC.t21 VCC.n82 0.814017
R1217 VCC.t15 VCC.n31 0.814017
R1218 VCC.n35 VCC.t15 0.814017
R1219 VCC.n222 VCC 0.799426
R1220 VCC.n151 VCC.n150 0.677583
R1221 VCC.n65 VCC.n64 0.6205
R1222 VCC.n66 VCC.n65 0.510369
R1223 VCC.n53 VCC.n52 0.490955
R1224 VCC VCC.n0 0.481269
R1225 VCC.n120 VCC.n119 0.434875
R1226 VCC.n105 VCC.n12 0.429597
R1227 VCC.n71 VCC.n66 0.423227
R1228 VCC.n97 VCC.n96 0.423227
R1229 VCC VCC.n148 0.335685
R1230 VCC.n94 VCC.n66 0.321523
R1231 VCC.n0 VCC 0.303385
R1232 VCC.n150 VCC.n149 0.298417
R1233 VCC VCC.n206 0.284691
R1234 VCC.n93 VCC.n92 0.280262
R1235 VCC.n134 VCC.n119 0.242167
R1236 VCC.n94 VCC.n93 0.224184
R1237 VCC.n149 VCC.n134 0.213463
R1238 VCC.n166 VCC 0.207566
R1239 VCC.n150 VCC.n119 0.161958
R1240 VCC.n92 VCC.n91 0.140381
R1241 VCC.n96 VCC 0.133783
R1242 VCC.n223 VCC.n105 0.128
R1243 VCC.n207 VCC 0.124875
R1244 VCC.n135 VCC 0.124875
R1245 VCC.n207 VCC 0.109601
R1246 VCC.n135 VCC 0.109601
R1247 VCC.n206 VCC.n205 0.108833
R1248 VCC.n219 VCC.n207 0.107956
R1249 VCC.n136 VCC.n135 0.105215
R1250 VCC.n134 VCC 0.0977222
R1251 VCC VCC.n165 0.0961731
R1252 VCC VCC.n0 0.0946265
R1253 VCC.n95 VCC.n94 0.0916778
R1254 VCC.n179 VCC.n166 0.0883378
R1255 VCC.n165 VCC 0.0868715
R1256 VCC.n165 VCC.n164 0.0855694
R1257 VCC.n95 VCC 0.0782027
R1258 VCC.n191 VCC.n181 0.0638663
R1259 VCC.n204 VCC.n194 0.0638663
R1260 VCC.n132 VCC.n121 0.0638663
R1261 VCC.n117 VCC.n116 0.0638663
R1262 VCC.n178 VCC.n167 0.0638663
R1263 VCC VCC.n133 0.0537407
R1264 VCC.n149 VCC 0.0525833
R1265 VCC VCC.n192 0.0484167
R1266 VCC.n205 VCC 0.0484167
R1267 VCC.n133 VCC.n120 0.0421667
R1268 VCC VCC.n223 0.0419157
R1269 VCC VCC.n179 0.0393514
R1270 VCC.n118 VCC 0.0359167
R1271 VCC.n93 VCC.n79 0.0268158
R1272 VCC.n96 VCC.n0 0.0178193
R1273 VCC.n149 VCC 0.00975926
R1274 VCC.n148 VCC.n136 0.00281481
R1275 VCC.n220 VCC.n219 0.00269298
R1276 VCC.n164 VCC.n152 0.00223611
R1277 VCC.n65 VCC.n53 0.00130906
R1278 COMPOUT.n2 COMPOUT.t2 113.796
R1279 COMPOUT.n6 COMPOUT.t3 84.6387
R1280 COMPOUT.n3 COMPOUT.t4 61.3556
R1281 COMPOUT.n5 COMPOUT.t0 41.6943
R1282 COMPOUT COMPOUT.t1 41.5734
R1283 COMPOUT.n7 COMPOUT.n6 3.52161
R1284 COMPOUT.n8 COMPOUT.n7 3.49783
R1285 COMPOUT.n7 COMPOUT.n2 2.22055
R1286 COMPOUT.n6 COMPOUT.n5 1.59772
R1287 COMPOUT.n8 COMPOUT 0.453774
R1288 COMPOUT.n5 COMPOUT.n4 0.323684
R1289 COMPOUT.n0 COMPOUT 0.208833
R1290 COMPOUT.n0 COMPOUT 0.179071
R1291 COMPOUT.n3 COMPOUT 0.119281
R1292 COMPOUT.n1 COMPOUT 0.0772045
R1293 COMPOUT.n1 COMPOUT.n0 0.0734167
R1294 COMPOUT COMPOUT.n8 0.0600238
R1295 COMPOUT.n4 COMPOUT 0.0587461
R1296 COMPOUT.n2 COMPOUT.n1 0.03225
R1297 COMPOUT.n4 COMPOUT.n3 0.0070445
R1298 x1.x2.x2.Z x1.x2.OUT.t1 113.781
R1299 x1.x1.ADJ x1.x2.OUT.t4 60.56
R1300 x1.x1.ADJ x1.x2.OUT.t3 53.3636
R1301 x1.x2.x2.Z x1.x2.OUT.t0 41.6352
R1302 x1.x2.x2.Z x1.x1.ADJ 6.3988
R1303 x1.x2.x2.Z x1.x2.OUT.t2 1.35076
R1304 CAL.n1 CAL.t6 234.692
R1305 CAL CAL.t0 233.88
R1306 CAL.n2 CAL.t5 229.185
R1307 CAL.n7 CAL.t1 193.226
R1308 CAL.n0 CAL.t3 193.153
R1309 CAL.n0 CAL.t2 174.048
R1310 CAL.n8 CAL.t4 174.005
R1311 CAL.n12 CAL.n0 12.9781
R1312 CAL.n1 CAL 4.63738
R1313 CAL.n3 CAL.n2 4.5005
R1314 CAL.n0 CAL 1.89741
R1315 CAL.n11 CAL.n10 1.46824
R1316 CAL.n7 CAL 1.188
R1317 CAL.n0 CAL 1.188
R1318 CAL.n10 CAL.n9 1.10352
R1319 CAL.n9 CAL.n6 1.09448
R1320 CAL.n3 CAL 1.04576
R1321 CAL.n9 CAL.n8 0.853
R1322 CAL.n13 CAL 0.721967
R1323 CAL.n13 CAL 0.6255
R1324 CAL.n6 CAL.n5 0.559652
R1325 CAL.n12 CAL.n11 0.203625
R1326 CAL.n5 CAL.n4 0.188
R1327 CAL.n4 CAL 0.180647
R1328 CAL.n6 CAL.n2 0.124054
R1329 CAL.n8 CAL.n7 0.0820074
R1330 CAL CAL.n12 0.063
R1331 CAL CAL.n13 0.0565538
R1332 CAL.n11 CAL 0.041125
R1333 CAL.n10 CAL.n1 0.0394785
R1334 CAL.n5 CAL 0.0194732
R1335 CAL.n4 CAL.n3 0.00481034
R1336 x1.x3.x2.GP x1.x3.SEL_N.t2 239.171
R1337 x1.x3.x3.GN x1.x3.SEL_N.t3 233.901
R1338 x1.x3.x2.GP x1.x3.SEL_N.t0 113.802
R1339 x1.x3.x2.GP x1.x3.SEL_N.t1 83.8505
R1340 x1.x3.x2.GP x1.x3.x3.GN 6.46588
R1341 EN_N.n3 EN_N.t0 1043.05
R1342 EN_N.t0 EN_N.n0 1040.82
R1343 EN_N.n0 EN_N.t2 194.654
R1344 EN_N.n2 EN_N.t3 7.78263
R1345 EN_N.n1 EN_N.t1 6.12265
R1346 EN_N.n2 EN_N.n1 2.50721
R1347 EN_N.n3 EN_N.n2 1.70148
R1348 EN_N.n5 EN_N.n4 1.66176
R1349 EN_N.n1 EN_N 1.2505
R1350 EN_N.n6 EN_N 1.2505
R1351 EN_N.n4 EN_N.n3 0.557375
R1352 EN_N.n5 EN_N 0.45675
R1353 EN_N.n4 EN_N.n0 0.163
R1354 EN_N.n1 EN_N 0.063
R1355 EN_N.n6 EN_N.n5 0.0510952
R1356 EN_N EN_N.n6 0.00645238
R1357 USEEXT.n0 USEEXT.t3 234.597
R1358 USEEXT.n1 USEEXT.t1 229.232
R1359 USEEXT.n5 USEEXT.t2 193.243
R1360 USEEXT.n6 USEEXT.t0 174.012
R1361 USEEXT.n0 USEEXT 4.63738
R1362 USEEXT.n2 USEEXT.n1 4.52679
R1363 USEEXT.n9 USEEXT.n8 1.313
R1364 USEEXT.n5 USEEXT 1.188
R1365 USEEXT.n8 USEEXT.n7 1.10352
R1366 USEEXT.n7 USEEXT.n4 1.09548
R1367 USEEXT.n7 USEEXT.n6 0.853
R1368 USEEXT.n4 USEEXT.n3 0.5005
R1369 USEEXT USEEXT.n9 0.195473
R1370 USEEXT.n10 USEEXT 0.129484
R1371 USEEXT.n4 USEEXT.n1 0.123161
R1372 USEEXT.n2 USEEXT 0.10425
R1373 USEEXT.n10 USEEXT 0.099413
R1374 USEEXT.n6 USEEXT.n5 0.0820074
R1375 USEEXT.n3 USEEXT.n2 0.0596518
R1376 USEEXT.n9 USEEXT 0.041125
R1377 USEEXT.n3 USEEXT 0.0339821
R1378 USEEXT USEEXT.n10 0.0236481
R1379 USEEXT.n8 USEEXT.n0 0.0218235
R1380 x3.x2.GP x3.SEL_N.t2 239.28
R1381 x3.x3.GN x3.SEL_N.t3 233.856
R1382 x3.x2.GP x3.SEL_N.t0 113.802
R1383 x3.x2.GP x3.SEL_N.t1 83.8505
R1384 x3.x2.GP x3.x3.GN 6.32014
R1385 x1.x3.OUT x1.x3.OUT.t1 113.803
R1386 x1.x3.OUT x1.x3.OUT.t2 113.796
R1387 x1.x3.OUT x1.x3.OUT.t4 68.4234
R1388 x1.x3.OUT x1.x3.OUT.t0 41.6342
R1389 x1.x3.OUT x1.x3.OUT.t3 41.507
R1390 x1.x3.OUT x1.x3.OUT.n0 7.4523
R1391 x1.x3.OUT.n0 x1.x3.OUT 2.78298
R1392 x1.x3.OUT.n0 x1.x3.OUT 1.90525
R1393 x1.x3.OUT.n0 x1.x3.OUT 1.89141
R1394 x3.OUT x3.OUT.t2 113.796
R1395 x3.OUT x3.OUT.t5 113.788
R1396 x3.OUT x3.OUT.t3 113.746
R1397 x3.OUT x3.OUT.t6 68.4093
R1398 x3.OUT x3.OUT.t4 41.6342
R1399 x3.OUT x3.OUT.t0 41.5734
R1400 x3.OUT x3.OUT.t1 41.4179
R1401 x3.OUT.n0 x3.OUT 7.4537
R1402 x3.OUT.n0 x3.OUT 1.81143
R1403 x3.OUT x3.OUT.n0 1.03936
R1404 x1.x1.inhigh x1.x1.inhigh.t2 115.745
R1405 x1.x1.inhigh x1.x1.inhigh.t1 31.1787
R1406 x1.x1.inhigh x1.x1.inhigh.t0 29.4286
R1407 DACOUT.n1 DACOUT.t2 113.761
R1408 DACOUT.n0 DACOUT.t1 41.6303
R1409 DACOUT DACOUT.n1 0.272792
R1410 DACOUT.n0 DACOUT 0.08175
R1411 DACOUT DACOUT.n0 0.0573182
R1412 DACOUT.n1 DACOUT 0.0402727
R1413 EXTTHRESH.n1 EXTTHRESH.t0 113.788
R1414 EXTTHRESH EXTTHRESH.t1 41.5734
R1415 EXTTHRESH.n2 EXTTHRESH.n1 8.40727
R1416 EXTTHRESH.n2 EXTTHRESH 0.39673
R1417 EXTTHRESH.n0 EXTTHRESH 0.08175
R1418 EXTTHRESH.n0 EXTTHRESH 0.0573182
R1419 EXTTHRESH EXTTHRESH.n2 0.0536915
R1420 EXTTHRESH.n1 EXTTHRESH.n0 0.0175455
R1421 INPUT.n1 INPUT.t0 113.761
R1422 INPUT INPUT.t1 41.5734
R1423 INPUT.n2 INPUT 1.2505
R1424 INPUT.n2 INPUT 0.70122
R1425 INPUT INPUT.n1 0.272792
R1426 INPUT.n1 INPUT.n0 0.0970909
R1427 INPUT.n0 INPUT 0.08175
R1428 INPUT.n0 INPUT 0.0573182
R1429 INPUT INPUT.n2 0.0421667
C0 VCC x1.x1.mirhigh 3.92074f
C1 x3.OUT x1.x3.OUT 1.39678f
C2 x1.x1.mirhigh COMPOUT 0.15303f
C3 CAL USEEXT 0.184631f
C4 VCC CAL 5.530931f
C5 x1.x1.mirhigh EN_N 0.736523f
C6 VCC USEEXT 2.91144f
C7 x1.x2.x2.GP CAL 1.13808f
C8 COMPOUT CAL 0.472262f
C9 x1.x1.mirhigh x1.x1.G1 0.00484f
C10 x1.x1.pg2g x1.x3.OUT 4.49e-19
C11 x1.x1.mirhigh x1.x1.G2 0.001507f
C12 x1.x3.OUT INPUT 0.624154f
C13 b6 b7 0.098267f
C14 VCC x1.x2.x2.GP 1.36206f
C15 VCC COMPOUT 1.97873f
C16 x1.x1.mirhigh x1.x1.inhigh 0.01694f
C17 VCC EN_N 11.370099f
C18 x1.x2.x2.GP COMPOUT 0.976261f
C19 CAL x1.x1.G1 0.026807f
C20 CAL x1.x1.G2 0.027326f
C21 EN_N COMPOUT 0.916628f
C22 VCC x1.x1.G1 1.49989f
C23 VCC x1.x1.G2 0.932067f
C24 b4 b3 0.098267f
C25 COMPOUT x1.x1.G1 0.010549f
C26 COMPOUT x1.x1.G2 0.471118f
C27 VCC x1.x1.inhigh 2.00666f
C28 EN_N x1.x1.G1 0.15289f
C29 EN_N x1.x1.G2 0.004728f
C30 x3.OUT INPUT 1.73035f
C31 USEEXT b7 0.095869f
C32 x3.OUT DACOUT 0.624154f
C33 a_9166_30798# DACOUT 0.106769f
C34 x1.x1.G1 x1.x1.G2 0.305193f
C35 EN_N x1.x1.inhigh 0.891479f
C36 a_7966_30798# a_7366_26366# 0.131455f
C37 VCC x1.x1.n2n 0.200319f
C38 x1.x1.mirhigh x1.x3.OUT 1.41e-19
C39 x1.x1.inhigh x1.x1.G1 0.896861f
C40 x1.x1.inhigh x1.x1.G2 0.104764f
C41 VCC x1.x1.p2p 0.888453f
C42 INPUT DACOUT 0.003124f
C43 x3.OUT EXTTHRESH 1.20931f
C44 b2 b3 0.098267f
C45 x1.x1.n2n EN_N 0.001021f
C46 CAL x1.x3.OUT 1.35366f
C47 a_6766_30798# a_7366_26366# 0.209322f
C48 VCC x1.x3.OUT 2.84465f
C49 x1.x1.n2n x1.x1.G1 0.676922f
C50 x1.x1.p2p EN_N 0.150607f
C51 b4 b5 0.098267f
C52 EXTTHRESH INPUT 0.068825f
C53 x1.x1.p2p x1.x1.G1 0.02214f
C54 x1.x1.n2n x1.x1.inhigh 5.52e-19
C55 EXTTHRESH DACOUT 0.47814f
C56 EN_N x1.x3.OUT 0.040617f
C57 b6 b5 0.098267f
C58 x1.x3.OUT x1.x1.G1 0.410051f
C59 x1.x3.OUT x1.x1.G2 1.28923f
C60 x3.OUT CAL 2.16026f
C61 x1.x1.mirhigh x1.x1.pg2g 1.02871f
C62 x3.OUT USEEXT 0.76179f
C63 a_9166_30798# USEEXT 4.46e-21
C64 x1.x1.inhigh x1.x3.OUT 0.692478f
C65 VCC x3.OUT 3.88477f
C66 a_6766_30798# a_5366_34798# 1.8e-21
C67 CAL INPUT 1.08969f
C68 USEEXT INPUT 0.054487f
C69 x3.OUT EN_N 0.235529f
C70 a_6166_26366# a_7366_26366# 0.182372f
C71 VCC x1.x1.pg2g 3.78855f
C72 a_6766_30798# a_6166_26366# 0.131455f
C73 VCC INPUT 0.349577f
C74 USEEXT DACOUT 1.0509f
C75 VCC DACOUT 0.301947f
C76 x3.OUT x1.x1.G1 1.40388f
C77 COMPOUT x1.x1.pg2g 1.16101f
C78 x3.OUT x1.x1.G2 0.036113f
C79 EN_N x1.x1.pg2g 0.022954f
C80 x3.OUT x1.x1.inhigh 0.729549f
C81 a_8566_26366# a_9166_30798# 0.131485f
C82 USEEXT EXTTHRESH 0.58553f
C83 x1.x1.pg2g x1.x1.G1 0.397601f
C84 a_7966_30798# a_8566_26366# 0.209322f
C85 x1.x1.pg2g x1.x1.G2 0.153401f
C86 b6 USEEXT 4.46e-21
C87 VCC EXTTHRESH 0.322957f
C88 x1.x1.inhigh x1.x1.pg2g 0.00845f
C89 x1.x1.n2n x3.OUT 0.001596f
C90 b1 b2 0.098267f
C91 a_5366_34798# a_6166_26366# 0.20932f
C92 b0 b1 0.098267f
C93 a_8566_26366# DACOUT 0.151801f
C94 a_8566_26366# a_7366_26366# 0.182372f
C95 USEEXT VSS 12.287024f
C96 EXTTHRESH VSS 2.741214f
C97 INPUT VSS 5.94419f
C98 CAL VSS 15.940003f
C99 COMPOUT VSS 7.38893f
C100 EN_N VSS 8.746689f
C101 DACOUT VSS 5.86254f
C102 b7 VSS 1.03263f
C103 b6 VSS 1.04109f
C104 b5 VSS 1.04109f
C105 b4 VSS 1.04109f
C106 b3 VSS 1.04109f
C107 b2 VSS 1.04109f
C108 b1 VSS 1.0411f
C109 b0 VSS 1.15272f
C110 VCC VSS 81.67105f
C111 x1.x2.x2.GP VSS 0.942725f
C112 x1.x1.pg2g VSS 4.93169f
C113 x1.x1.G2 VSS 9.06897f
C114 x1.x3.OUT VSS 6.916137f
C115 x3.OUT VSS 17.223436f
C116 x1.x1.n2n VSS 0.996702f
C117 x1.x1.G1 VSS 7.98487f
C118 x1.x1.mirhigh VSS 1.527153f
C119 x1.x1.inhigh VSS 2.94796f
C120 x1.x1.p2p VSS 0.150606f
C121 a_9166_30798# VSS 2.28437f
C122 a_8566_26366# VSS 6.30451f
C123 a_7966_30798# VSS 2.2293f
C124 a_7366_26366# VSS 6.29855f
C125 a_6766_30798# VSS 2.23322f
C126 a_6166_26366# VSS 6.44599f
C127 a_5366_34798# VSS 5.98194f
C128 EXTTHRESH.t0 VSS 0.033179f
C129 EXTTHRESH.t1 VSS 0.032061f
C130 EXTTHRESH.n0 VSS 0.042376f
C131 EXTTHRESH.n1 VSS 0.814215f
C132 EXTTHRESH.n2 VSS 0.690785f
C133 x1.x1.inhigh.t2 VSS 0.040812f
C134 x1.x1.inhigh.t1 VSS 0.141031f
C135 x1.x1.inhigh.t0 VSS 0.141031f
C136 x3.OUT.t5 VSS 0.023972f
C137 x3.OUT.t1 VSS 0.022658f
C138 x3.OUT.t3 VSS 0.02392f
C139 x3.OUT.t2 VSS 0.023987f
C140 x3.OUT.t4 VSS 0.023227f
C141 x3.OUT.n0 VSS 0.786911f
C142 x3.OUT.t6 VSS 0.489025f
C143 x3.OUT.t0 VSS 0.023165f
C144 x1.x3.OUT.n0 VSS 1.19689f
C145 x1.x3.OUT.t2 VSS 0.014249f
C146 x1.x3.OUT.t4 VSS 0.290549f
C147 x1.x3.OUT.t3 VSS 0.013538f
C148 x1.x3.OUT.t1 VSS 0.014256f
C149 x1.x3.OUT.t0 VSS 0.013797f
C150 x3.x2.GP VSS 1.21235f
C151 x3.SEL_N.t2 VSS 0.023121f
C152 x3.SEL_N.t3 VSS 0.02306f
C153 x3.x3.GN VSS 0.8024f
C154 x3.SEL_N.t1 VSS 0.01268f
C155 x3.SEL_N.t0 VSS 0.026393f
C156 USEEXT.t3 VSS 0.009857f
C157 USEEXT.n0 VSS 0.066754f
C158 USEEXT.t1 VSS 0.009705f
C159 USEEXT.n1 VSS 0.07375f
C160 USEEXT.n2 VSS 0.02639f
C161 USEEXT.n3 VSS 0.011056f
C162 USEEXT.n4 VSS 0.052399f
C163 USEEXT.t2 VSS 0.005772f
C164 USEEXT.n5 VSS 0.082707f
C165 USEEXT.t0 VSS 0.017774f
C166 USEEXT.n6 VSS 0.080674f
C167 USEEXT.n7 VSS 0.249377f
C168 USEEXT.n8 VSS 0.052528f
C169 USEEXT.n9 VSS 0.029834f
C170 USEEXT.n10 VSS 0.033799f
C171 EN_N.t2 VSS 0.043622f
C172 EN_N.n0 VSS 2.33303f
C173 EN_N.t1 VSS 1.25083f
C174 EN_N.n1 VSS 1.50456f
C175 EN_N.t3 VSS 1.7794f
C176 EN_N.n2 VSS 2.31188f
C177 EN_N.t0 VSS 0.052172f
C178 EN_N.n3 VSS 0.949479f
C179 EN_N.n4 VSS 0.563693f
C180 EN_N.n5 VSS 0.266324f
C181 EN_N.n6 VSS 0.029419f
C182 x1.x3.x2.GP VSS 1.20755f
C183 x1.x3.SEL_N.t2 VSS 0.023118f
C184 x1.x3.SEL_N.t3 VSS 0.023076f
C185 x1.x3.x3.GN VSS 0.807187f
C186 x1.x3.SEL_N.t0 VSS 0.026392f
C187 x1.x3.SEL_N.t1 VSS 0.01268f
C188 CAL.t3 VSS 0.013208f
C189 CAL.t2 VSS 0.04076f
C190 CAL.t0 VSS 0.025293f
C191 CAL.n0 VSS 1.68117f
C192 CAL.t6 VSS 0.022602f
C193 CAL.n1 VSS 0.141658f
C194 CAL.t5 VSS 0.022188f
C195 CAL.n2 VSS 0.168561f
C196 CAL.n3 VSS 0.005959f
C197 CAL.n4 VSS 0.008409f
C198 CAL.n5 VSS 0.070479f
C199 CAL.n6 VSS 0.125859f
C200 CAL.t4 VSS 0.040717f
C201 CAL.t1 VSS 0.01327f
C202 CAL.n7 VSS 0.194094f
C203 CAL.n8 VSS 0.187827f
C204 CAL.n9 VSS 0.569952f
C205 CAL.n10 VSS 0.039611f
C206 CAL.n11 VSS 0.054454f
C207 CAL.n12 VSS 0.754326f
C208 CAL.n13 VSS 0.142505f
C209 x1.x2.OUT.t2 VSS 1.20129f
C210 x1.x2.x2.Z VSS 0.787408f
C211 x1.x1.ADJ VSS 0.102848f
C212 x1.x2.OUT.t3 VSS 0.002626f
C213 x1.x2.OUT.t4 VSS 0.003534f
C214 x1.x2.OUT.t1 VSS 0.001163f
C215 x1.x2.OUT.t0 VSS 0.001127f
C216 VCC.n0 VSS 0.567249f
C217 VCC.t22 VSS 0.570362f
C218 VCC.n1 VSS 0.018498f
C219 VCC.n2 VSS 0.018582f
C220 VCC.n4 VSS 0.018923f
C221 VCC.n5 VSS 0.018907f
C222 VCC.n6 VSS 0.131033f
C223 VCC.t13 VSS 0.188556f
C224 VCC.n8 VSS 0.018923f
C225 VCC.n9 VSS 0.131033f
C226 VCC.n10 VSS 0.013263f
C227 VCC.n11 VSS 0.013229f
C228 VCC.n12 VSS 0.587609f
C229 VCC.n13 VSS 0.0288f
C230 VCC.n14 VSS 0.023581f
C231 VCC.n15 VSS 0.403177f
C232 VCC.n16 VSS 0.403177f
C233 VCC.n17 VSS 0.027454f
C234 VCC.n18 VSS 0.039177f
C235 VCC.n19 VSS 0.039988f
C236 VCC.n21 VSS 0.041215f
C237 VCC.n22 VSS 0.041208f
C238 VCC.n23 VSS 0.466789f
C239 VCC.t17 VSS 0.761721f
C240 VCC.n25 VSS 0.041215f
C241 VCC.n26 VSS 0.466789f
C242 VCC.n27 VSS 0.033749f
C243 VCC.n28 VSS 0.034039f
C244 VCC.n29 VSS 0.037772f
C245 VCC.n30 VSS 0.04894f
C246 VCC.n32 VSS 0.04894f
C247 VCC.n33 VSS 0.048347f
C248 VCC.n34 VSS 0.527106f
C249 VCC.t15 VSS 0.806632f
C250 VCC.n36 VSS 0.04894f
C251 VCC.n37 VSS 0.527106f
C252 VCC.n38 VSS 0.034241f
C253 VCC.n39 VSS 0.041164f
C254 VCC.n40 VSS 0.458848f
C255 VCC.n41 VSS 0.025251f
C256 VCC.n42 VSS 0.041215f
C257 VCC.n43 VSS 0.041215f
C258 VCC.t16 VSS 0.761721f
C259 VCC.n44 VSS 0.040355f
C260 VCC.n46 VSS 0.466789f
C261 VCC.n47 VSS 0.041215f
C262 VCC.n49 VSS 0.466789f
C263 VCC.n50 VSS 0.040228f
C264 VCC.n51 VSS 0.028004f
C265 VCC.n52 VSS 1.31232f
C266 VCC.t19 VSS 0.058269f
C267 VCC.n53 VSS 0.722939f
C268 VCC.n54 VSS 0.028563f
C269 VCC.n55 VSS 0.03021f
C270 VCC.n56 VSS 0.03021f
C271 VCC.t18 VSS 0.327871f
C272 VCC.n57 VSS 0.033078f
C273 VCC.n59 VSS 0.198721f
C274 VCC.n60 VSS 0.03021f
C275 VCC.n62 VSS 0.198721f
C276 VCC.n63 VSS 0.033132f
C277 VCC.n64 VSS 0.028474f
C278 VCC.n65 VSS 0.554276f
C279 VCC.n66 VSS 0.71706f
C280 VCC.t3 VSS 0.023237f
C281 VCC.n67 VSS 0.028204f
C282 VCC.n68 VSS 0.050703f
C283 VCC.n69 VSS 0.519154f
C284 VCC.n70 VSS 0.519154f
C285 VCC.n71 VSS 0.046745f
C286 VCC.n72 VSS 0.046827f
C287 VCC.n73 VSS 0.048353f
C288 VCC.t2 VSS 0.884041f
C289 VCC.n76 VSS 0.048353f
C290 VCC.n77 VSS 0.047512f
C291 VCC.n78 VSS 0.026695f
C292 VCC.n79 VSS 0.049749f
C293 VCC.n80 VSS 0.034279f
C294 VCC.n81 VSS 0.04894f
C295 VCC.n83 VSS 0.04894f
C296 VCC.n84 VSS 0.048347f
C297 VCC.n85 VSS 0.527106f
C298 VCC.t21 VSS 0.806632f
C299 VCC.n87 VSS 0.04894f
C300 VCC.n88 VSS 0.527106f
C301 VCC.n89 VSS 0.037572f
C302 VCC.n90 VSS 0.047789f
C303 VCC.t12 VSS 0.011655f
C304 VCC.n91 VSS 0.0701f
C305 VCC.n92 VSS 0.265565f
C306 VCC.n93 VSS 0.062721f
C307 VCC.n94 VSS 0.390108f
C308 VCC.n95 VSS 0.045082f
C309 VCC.n96 VSS 0.45358f
C310 VCC.n97 VSS 0.050728f
C311 VCC.n98 VSS 0.051196f
C312 VCC.n99 VSS 0.04456f
C313 VCC.t11 VSS 0.673282f
C314 VCC.n102 VSS 0.04456f
C315 VCC.n103 VSS 0.043878f
C316 VCC.n104 VSS 0.024328f
C317 VCC.n105 VSS 0.156637f
C318 VCC.n106 VSS 0.01622f
C319 VCC.n107 VSS 0.067835f
C320 VCC.n108 VSS 0.019387f
C321 VCC.n109 VSS 0.019387f
C322 VCC.n110 VSS 0.013746f
C323 VCC.n111 VSS 0.01993f
C324 VCC.n112 VSS 0.119873f
C325 VCC.t14 VSS 0.195783f
C326 VCC.n115 VSS 0.119873f
C327 VCC.n116 VSS 0.044082f
C328 VCC.n117 VSS 0.01853f
C329 VCC.n118 VSS 0.29565f
C330 VCC.n119 VSS 0.348745f
C331 VCC.n120 VSS 0.288015f
C332 VCC.n121 VSS 0.044082f
C333 VCC.n122 VSS 0.019888f
C334 VCC.n123 VSS 0.019888f
C335 VCC.n124 VSS 0.019888f
C336 VCC.n125 VSS 0.070724f
C337 VCC.n126 VSS 0.013767f
C338 VCC.n127 VSS 0.128916f
C339 VCC.t5 VSS 0.176696f
C340 VCC.n130 VSS 0.128916f
C341 VCC.n131 VSS 0.016241f
C342 VCC.n132 VSS 0.01853f
C343 VCC.n133 VSS 0.030248f
C344 VCC.n134 VSS 0.193947f
C345 VCC.n135 VSS 0.070343f
C346 VCC.t8 VSS 0.023222f
C347 VCC.n136 VSS 0.060251f
C348 VCC.n137 VSS 0.013813f
C349 VCC.n138 VSS 0.01997f
C350 VCC.n139 VSS 0.01997f
C351 VCC.t7 VSS 0.202862f
C352 VCC.n140 VSS 0.020082f
C353 VCC.n142 VSS 0.130604f
C354 VCC.n143 VSS 0.01997f
C355 VCC.n145 VSS 0.130604f
C356 VCC.n146 VSS 0.020024f
C357 VCC.n147 VSS 0.013792f
C358 VCC.n148 VSS 0.107568f
C359 VCC.n149 VSS 0.208538f
C360 VCC.n150 VSS 0.367728f
C361 VCC.n151 VSS 0.551199f
C362 VCC.t1 VSS 0.023215f
C363 VCC.n152 VSS 0.271819f
C364 VCC.n153 VSS 0.013813f
C365 VCC.n154 VSS 0.01997f
C366 VCC.n155 VSS 0.01997f
C367 VCC.t0 VSS 0.202862f
C368 VCC.n156 VSS 0.020082f
C369 VCC.n158 VSS 0.130604f
C370 VCC.n159 VSS 0.01997f
C371 VCC.n161 VSS 0.130604f
C372 VCC.n162 VSS 0.020024f
C373 VCC.n163 VSS 0.013792f
C374 VCC.n164 VSS 0.031477f
C375 VCC.n165 VSS 0.090443f
C376 VCC.n166 VSS 0.179951f
C377 VCC.n167 VSS 0.044082f
C378 VCC.n168 VSS 0.019888f
C379 VCC.n169 VSS 0.019888f
C380 VCC.n170 VSS 0.019888f
C381 VCC.n171 VSS 0.066908f
C382 VCC.n172 VSS 0.013767f
C383 VCC.n173 VSS 0.128916f
C384 VCC.t20 VSS 0.176696f
C385 VCC.n176 VSS 0.128916f
C386 VCC.n177 VSS 0.016241f
C387 VCC.n178 VSS 0.01853f
C388 VCC.n179 VSS 0.075824f
C389 VCC.n180 VSS 0.068439f
C390 VCC.n181 VSS 0.044082f
C391 VCC.n182 VSS 0.019888f
C392 VCC.n183 VSS 0.019888f
C393 VCC.n184 VSS 0.019888f
C394 VCC.n185 VSS 0.013767f
C395 VCC.n186 VSS 0.128916f
C396 VCC.t4 VSS 0.176696f
C397 VCC.n189 VSS 0.128916f
C398 VCC.n190 VSS 0.016241f
C399 VCC.n191 VSS 0.01853f
C400 VCC.n192 VSS 0.193934f
C401 VCC.n193 VSS 0.066908f
C402 VCC.n194 VSS 0.044082f
C403 VCC.n195 VSS 0.01993f
C404 VCC.n196 VSS 0.119873f
C405 VCC.n197 VSS 0.119873f
C406 VCC.n198 VSS 0.013746f
C407 VCC.n199 VSS 0.019387f
C408 VCC.t6 VSS 0.195783f
C409 VCC.n202 VSS 0.019387f
C410 VCC.n203 VSS 0.01622f
C411 VCC.n204 VSS 0.01853f
C412 VCC.n205 VSS 0.061479f
C413 VCC.n206 VSS 0.152704f
C414 VCC.n207 VSS 0.070966f
C415 VCC.n208 VSS 0.013836f
C416 VCC.n209 VSS 0.02001f
C417 VCC.n210 VSS 0.136697f
C418 VCC.n211 VSS 0.136697f
C419 VCC.n212 VSS 0.020039f
C420 VCC.n213 VSS 0.020421f
C421 VCC.t9 VSS 0.189775f
C422 VCC.n216 VSS 0.020421f
C423 VCC.n217 VSS 0.019981f
C424 VCC.n218 VSS 0.013816f
C425 VCC.n219 VSS 0.02492f
C426 VCC.t10 VSS 0.023215f
C427 VCC.n220 VSS 0.214959f
C428 VCC.n221 VSS 1.45106f
C429 VCC.n222 VSS 2.71235f
C430 VCC.n223 VSS 1.26026f
C431 x1.x1.mirhigh.t1 VSS 0.241652f
C432 x1.x1.mirhigh.t0 VSS 0.472059f
C433 x1.x1.mirhigh.t2 VSS 0.294208f
C434 x1.x1.mirhigh.n0 VSS 2.23501f
C435 x1.x1.pg2g.t2 VSS 0.771449f
C436 x1.x1.pg2g.t0 VSS 0.738093f
C437 x1.x1.pg2g.t1 VSS 0.060558f
.ends

