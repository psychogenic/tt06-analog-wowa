magic
tech sky130A
magscale 1 2
timestamp 1713327229
<< viali >>
rect 1409 14569 1443 14603
rect 2053 14569 2087 14603
rect 3065 14569 3099 14603
rect 4077 14569 4111 14603
rect 5089 14569 5123 14603
rect 6377 14569 6411 14603
rect 7113 14569 7147 14603
rect 8125 14569 8159 14603
rect 9137 14569 9171 14603
rect 13369 14501 13403 14535
rect 1593 14365 1627 14399
rect 2237 14365 2271 14399
rect 3249 14365 3283 14399
rect 4261 14365 4295 14399
rect 5273 14365 5307 14399
rect 6561 14365 6595 14399
rect 7297 14365 7331 14399
rect 8309 14365 8343 14399
rect 9321 14365 9355 14399
rect 11161 14365 11195 14399
rect 12357 14365 12391 14399
rect 13185 14365 13219 14399
rect 11345 14229 11379 14263
rect 12173 14229 12207 14263
rect 3525 14025 3559 14059
rect 4537 14025 4571 14059
rect 3617 13957 3651 13991
rect 4169 13957 4203 13991
rect 7113 13957 7147 13991
rect 7297 13957 7331 13991
rect 3249 13889 3283 13923
rect 3709 13889 3743 13923
rect 3985 13889 4019 13923
rect 4261 13889 4295 13923
rect 4353 13889 4387 13923
rect 4629 13889 4663 13923
rect 6656 13911 6690 13945
rect 6929 13923 6963 13957
rect 6745 13889 6779 13923
rect 7021 13889 7055 13923
rect 9045 13889 9079 13923
rect 9229 13889 9263 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 10977 13889 11011 13923
rect 9137 13821 9171 13855
rect 4353 13753 4387 13787
rect 6929 13753 6963 13787
rect 3249 13685 3283 13719
rect 3341 13685 3375 13719
rect 3985 13685 4019 13719
rect 7297 13685 7331 13719
rect 10701 13685 10735 13719
rect 3433 13481 3467 13515
rect 5181 13481 5215 13515
rect 6193 13481 6227 13515
rect 6285 13481 6319 13515
rect 6837 13481 6871 13515
rect 2881 13413 2915 13447
rect 5549 13413 5583 13447
rect 3801 13345 3835 13379
rect 1501 13277 1535 13311
rect 3065 13277 3099 13311
rect 3525 13277 3559 13311
rect 5825 13277 5859 13311
rect 6285 13277 6319 13311
rect 6469 13277 6503 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 10066 13277 10100 13311
rect 10333 13277 10367 13311
rect 10425 13277 10459 13311
rect 1768 13209 1802 13243
rect 4046 13209 4080 13243
rect 5365 13209 5399 13243
rect 5917 13209 5951 13243
rect 6561 13209 6595 13243
rect 7450 13209 7484 13243
rect 10692 13209 10726 13243
rect 3157 13141 3191 13175
rect 3249 13141 3283 13175
rect 3525 13141 3559 13175
rect 6009 13141 6043 13175
rect 6653 13141 6687 13175
rect 6929 13141 6963 13175
rect 8585 13141 8619 13175
rect 8953 13141 8987 13175
rect 11805 13141 11839 13175
rect 2145 12937 2179 12971
rect 4629 12937 4663 12971
rect 4905 12937 4939 12971
rect 7941 12937 7975 12971
rect 9689 12937 9723 12971
rect 9873 12937 9907 12971
rect 11529 12937 11563 12971
rect 12173 12937 12207 12971
rect 5073 12869 5107 12903
rect 5273 12869 5307 12903
rect 12265 12869 12299 12903
rect 2329 12801 2363 12835
rect 3249 12801 3283 12835
rect 3505 12801 3539 12835
rect 6561 12801 6595 12835
rect 6817 12801 6851 12835
rect 9321 12801 9355 12835
rect 9870 12801 9904 12835
rect 10701 12801 10735 12835
rect 10885 12801 10919 12835
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 12541 12801 12575 12835
rect 9229 12733 9263 12767
rect 10333 12733 10367 12767
rect 11713 12733 11747 12767
rect 11805 12733 11839 12767
rect 12357 12733 12391 12767
rect 10793 12665 10827 12699
rect 5089 12597 5123 12631
rect 8953 12597 8987 12631
rect 9229 12597 9263 12631
rect 10241 12597 10275 12631
rect 10517 12597 10551 12631
rect 12357 12597 12391 12631
rect 12725 12597 12759 12631
rect 4813 12393 4847 12427
rect 5549 12393 5583 12427
rect 5733 12393 5767 12427
rect 5825 12393 5859 12427
rect 5987 12393 6021 12427
rect 6561 12393 6595 12427
rect 6745 12393 6779 12427
rect 9781 12393 9815 12427
rect 2237 12325 2271 12359
rect 9045 12325 9079 12359
rect 2973 12257 3007 12291
rect 11161 12257 11195 12291
rect 11529 12257 11563 12291
rect 11621 12257 11655 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 3157 12189 3191 12223
rect 5181 12189 5215 12223
rect 9229 12189 9263 12223
rect 9960 12189 9994 12223
rect 10277 12189 10311 12223
rect 10425 12189 10459 12223
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 10793 12189 10827 12223
rect 10885 12189 10919 12223
rect 11253 12189 11287 12223
rect 11437 12189 11471 12223
rect 11805 12189 11839 12223
rect 12081 12189 12115 12223
rect 12348 12189 12382 12223
rect 4767 12155 4801 12189
rect 2513 12121 2547 12155
rect 4997 12121 5031 12155
rect 6193 12121 6227 12155
rect 6377 12121 6411 12155
rect 10057 12121 10091 12155
rect 10149 12121 10183 12155
rect 2053 12053 2087 12087
rect 2697 12053 2731 12087
rect 4629 12053 4663 12087
rect 5549 12053 5583 12087
rect 5983 12053 6017 12087
rect 6587 12053 6621 12087
rect 9321 12053 9355 12087
rect 9413 12053 9447 12087
rect 9597 12053 9631 12087
rect 11989 12053 12023 12087
rect 13461 12053 13495 12087
rect 2973 11849 3007 11883
rect 3433 11849 3467 11883
rect 3709 11849 3743 11883
rect 4813 11849 4847 11883
rect 5089 11849 5123 11883
rect 5181 11849 5215 11883
rect 6377 11849 6411 11883
rect 7021 11849 7055 11883
rect 8493 11849 8527 11883
rect 10425 11849 10459 11883
rect 10793 11849 10827 11883
rect 11161 11849 11195 11883
rect 11621 11849 11655 11883
rect 12725 11849 12759 11883
rect 4721 11781 4755 11815
rect 4997 11781 5031 11815
rect 5733 11781 5767 11815
rect 6529 11781 6563 11815
rect 6745 11781 6779 11815
rect 7481 11781 7515 11815
rect 8033 11781 8067 11815
rect 9137 11781 9171 11815
rect 10241 11781 10275 11815
rect 12265 11781 12299 11815
rect 12357 11781 12391 11815
rect 4491 11747 4525 11781
rect 1501 11713 1535 11747
rect 1768 11713 1802 11747
rect 3157 11713 3191 11747
rect 3525 11713 3559 11747
rect 4077 11713 4111 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 7205 11713 7239 11747
rect 8677 11713 8711 11747
rect 9505 11713 9539 11747
rect 9689 11713 9723 11747
rect 10149 11713 10183 11747
rect 10333 11713 10367 11747
rect 10609 11713 10643 11747
rect 10701 11713 10735 11747
rect 10977 11713 11011 11747
rect 11253 11713 11287 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12081 11713 12115 11747
rect 12173 11713 12207 11747
rect 12541 11713 12575 11747
rect 13001 11713 13035 11747
rect 3249 11645 3283 11679
rect 3617 11645 3651 11679
rect 3893 11645 3927 11679
rect 3985 11645 4019 11679
rect 4169 11645 4203 11679
rect 5457 11645 5491 11679
rect 7297 11645 7331 11679
rect 8861 11645 8895 11679
rect 10425 11645 10459 11679
rect 12909 11645 12943 11679
rect 4353 11577 4387 11611
rect 5365 11577 5399 11611
rect 6009 11577 6043 11611
rect 7849 11577 7883 11611
rect 2881 11509 2915 11543
rect 4537 11509 4571 11543
rect 6561 11509 6595 11543
rect 7389 11509 7423 11543
rect 9045 11509 9079 11543
rect 9689 11509 9723 11543
rect 1685 11305 1719 11339
rect 2421 11305 2455 11339
rect 4445 11305 4479 11339
rect 6285 11305 6319 11339
rect 7113 11305 7147 11339
rect 7389 11305 7423 11339
rect 8401 11305 8435 11339
rect 12081 11305 12115 11339
rect 2237 11237 2271 11271
rect 7481 11237 7515 11271
rect 7941 11237 7975 11271
rect 8677 11237 8711 11271
rect 11529 11237 11563 11271
rect 12357 11237 12391 11271
rect 2697 11169 2731 11203
rect 3157 11169 3191 11203
rect 3801 11169 3835 11203
rect 4537 11169 4571 11203
rect 8217 11169 8251 11203
rect 10701 11169 10735 11203
rect 11897 11169 11931 11203
rect 1869 11101 1903 11135
rect 2789 11101 2823 11135
rect 2927 11101 2961 11135
rect 4077 11101 4111 11135
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 5273 11101 5307 11135
rect 5641 11101 5675 11135
rect 6377 11101 6411 11135
rect 6561 11101 6595 11135
rect 6653 11101 6687 11135
rect 6837 11101 6871 11135
rect 6929 11101 6963 11135
rect 7573 11101 7607 11135
rect 7849 11101 7883 11135
rect 8125 11101 8159 11135
rect 8493 11101 8527 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 10977 11101 11011 11135
rect 11253 11101 11287 11135
rect 11621 11101 11655 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 12081 11101 12115 11135
rect 12357 11101 12391 11135
rect 12633 11101 12667 11135
rect 13369 11101 13403 11135
rect 1961 11033 1995 11067
rect 2513 11033 2547 11067
rect 3065 11033 3099 11067
rect 4629 11033 4663 11067
rect 6126 11033 6160 11067
rect 8401 11033 8435 11067
rect 4169 10965 4203 10999
rect 4261 10965 4295 10999
rect 5917 10965 5951 10999
rect 6009 10965 6043 10999
rect 7757 10965 7791 10999
rect 12541 10965 12575 10999
rect 13185 10965 13219 10999
rect 3617 10761 3651 10795
rect 3899 10761 3933 10795
rect 4077 10761 4111 10795
rect 4445 10761 4479 10795
rect 4905 10761 4939 10795
rect 5457 10761 5491 10795
rect 7297 10761 7331 10795
rect 8585 10761 8619 10795
rect 11529 10761 11563 10795
rect 12633 10761 12667 10795
rect 6469 10693 6503 10727
rect 11687 10693 11721 10727
rect 11897 10693 11931 10727
rect 13369 10693 13403 10727
rect 3985 10625 4019 10659
rect 4721 10625 4755 10659
rect 4813 10625 4847 10659
rect 5733 10625 5767 10659
rect 6193 10625 6227 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 7142 10625 7176 10659
rect 7488 10625 7522 10659
rect 7757 10625 7791 10659
rect 8401 10625 8435 10659
rect 8769 10625 8803 10659
rect 8953 10625 8987 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 10701 10625 10735 10659
rect 10977 10625 11011 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 12265 10625 12299 10659
rect 12909 10625 12943 10659
rect 13553 10625 13587 10659
rect 4353 10557 4387 10591
rect 5181 10557 5215 10591
rect 6929 10557 6963 10591
rect 7573 10557 7607 10591
rect 13277 10557 13311 10591
rect 4261 10489 4295 10523
rect 5089 10489 5123 10523
rect 5917 10489 5951 10523
rect 9137 10489 9171 10523
rect 9597 10489 9631 10523
rect 10793 10489 10827 10523
rect 10885 10489 10919 10523
rect 11989 10489 12023 10523
rect 5825 10421 5859 10455
rect 6009 10421 6043 10455
rect 6745 10421 6779 10455
rect 7757 10421 7791 10455
rect 8769 10421 8803 10455
rect 9413 10421 9447 10455
rect 10057 10421 10091 10455
rect 10517 10421 10551 10455
rect 11713 10421 11747 10455
rect 4261 10217 4295 10251
rect 6653 10217 6687 10251
rect 7021 10217 7055 10251
rect 7665 10217 7699 10251
rect 7849 10217 7883 10251
rect 8953 10217 8987 10251
rect 11897 10217 11931 10251
rect 6193 10149 6227 10183
rect 6469 10149 6503 10183
rect 7481 10149 7515 10183
rect 12725 10149 12759 10183
rect 3893 10081 3927 10115
rect 7205 10081 7239 10115
rect 10333 10081 10367 10115
rect 4077 10013 4111 10047
rect 6561 10013 6595 10047
rect 6929 10013 6963 10047
rect 7021 10013 7055 10047
rect 7297 10013 7331 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 8585 10013 8619 10047
rect 12449 10013 12483 10047
rect 13093 10013 13127 10047
rect 6101 9945 6135 9979
rect 10066 9945 10100 9979
rect 10609 9945 10643 9979
rect 4629 9877 4663 9911
rect 6837 9877 6871 9911
rect 8677 9877 8711 9911
rect 5089 9673 5123 9707
rect 10057 9673 10091 9707
rect 10241 9673 10275 9707
rect 11897 9673 11931 9707
rect 6837 9605 6871 9639
rect 6929 9605 6963 9639
rect 11529 9605 11563 9639
rect 3249 9537 3283 9571
rect 5273 9537 5307 9571
rect 5549 9537 5583 9571
rect 6561 9537 6595 9571
rect 7113 9537 7147 9571
rect 7297 9537 7331 9571
rect 9045 9537 9079 9571
rect 9137 9537 9171 9571
rect 9413 9537 9447 9571
rect 9597 9537 9631 9571
rect 9689 9537 9723 9571
rect 9781 9537 9815 9571
rect 10149 9559 10183 9593
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11161 9537 11195 9571
rect 11713 9537 11747 9571
rect 12081 9537 12115 9571
rect 12337 9537 12371 9571
rect 2237 9469 2271 9503
rect 3065 9469 3099 9503
rect 3157 9469 3191 9503
rect 3341 9469 3375 9503
rect 5457 9469 5491 9503
rect 6745 9469 6779 9503
rect 9321 9469 9355 9503
rect 10885 9469 10919 9503
rect 10977 9469 11011 9503
rect 11345 9469 11379 9503
rect 2605 9401 2639 9435
rect 2881 9401 2915 9435
rect 9229 9401 9263 9435
rect 13461 9401 13495 9435
rect 2697 9333 2731 9367
rect 5549 9333 5583 9367
rect 6377 9333 6411 9367
rect 6837 9333 6871 9367
rect 10425 9333 10459 9367
rect 1501 9129 1535 9163
rect 2973 9129 3007 9163
rect 6745 9129 6779 9163
rect 9781 9129 9815 9163
rect 9965 9129 9999 9163
rect 11253 9129 11287 9163
rect 5089 9061 5123 9095
rect 3617 8993 3651 9027
rect 4813 8993 4847 9027
rect 5181 8993 5215 9027
rect 10057 8993 10091 9027
rect 11161 8993 11195 9027
rect 12081 8993 12115 9027
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3525 8925 3559 8959
rect 3985 8925 4019 8959
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 5917 8925 5951 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6837 8925 6871 8959
rect 9965 8925 9999 8959
rect 10425 8925 10459 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 10793 8925 10827 8959
rect 10977 8925 11011 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11805 8925 11839 8959
rect 11897 8925 11931 8959
rect 2614 8857 2648 8891
rect 10609 8857 10643 8891
rect 11621 8857 11655 8891
rect 12326 8857 12360 8891
rect 3341 8789 3375 8823
rect 3801 8789 3835 8823
rect 5549 8789 5583 8823
rect 6377 8789 6411 8823
rect 13461 8789 13495 8823
rect 1961 8585 1995 8619
rect 4169 8585 4203 8619
rect 4445 8585 4479 8619
rect 6193 8585 6227 8619
rect 6745 8585 6779 8619
rect 7389 8585 7423 8619
rect 7849 8585 7883 8619
rect 12173 8585 12207 8619
rect 12633 8585 12667 8619
rect 3740 8517 3774 8551
rect 4537 8517 4571 8551
rect 9321 8517 9355 8551
rect 2329 8449 2363 8483
rect 2421 8449 2455 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4629 8449 4663 8483
rect 5825 8449 5859 8483
rect 6469 8449 6503 8483
rect 6653 8449 6687 8483
rect 7205 8449 7239 8483
rect 7481 8449 7515 8483
rect 10149 8449 10183 8483
rect 10425 8449 10459 8483
rect 10793 8449 10827 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 12817 8449 12851 8483
rect 13001 8449 13035 8483
rect 2145 8381 2179 8415
rect 2237 8381 2271 8415
rect 5917 8381 5951 8415
rect 11069 8381 11103 8415
rect 2605 8313 2639 8347
rect 7021 8313 7055 8347
rect 4261 8245 4295 8279
rect 6009 8245 6043 8279
rect 6929 8245 6963 8279
rect 3341 8041 3375 8075
rect 5089 8041 5123 8075
rect 6377 8041 6411 8075
rect 6837 8041 6871 8075
rect 8217 8041 8251 8075
rect 8953 8041 8987 8075
rect 9597 8041 9631 8075
rect 10333 8041 10367 8075
rect 10701 8041 10735 8075
rect 3065 7973 3099 8007
rect 4997 7973 5031 8007
rect 9321 7973 9355 8007
rect 1685 7905 1719 7939
rect 6218 7905 6252 7939
rect 6561 7905 6595 7939
rect 6929 7905 6963 7939
rect 7021 7905 7055 7939
rect 9781 7894 9815 7928
rect 3525 7837 3559 7871
rect 3617 7837 3651 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5273 7837 5307 7871
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 5740 7837 5774 7871
rect 6009 7837 6043 7871
rect 7297 7837 7331 7871
rect 8493 7837 8527 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9505 7837 9539 7871
rect 10517 7837 10551 7871
rect 10793 7837 10827 7871
rect 1952 7769 1986 7803
rect 3341 7769 3375 7803
rect 6101 7701 6135 7735
rect 7205 7701 7239 7735
rect 8033 7701 8067 7735
rect 9781 7701 9815 7735
rect 5549 7497 5583 7531
rect 6653 7497 6687 7531
rect 7573 7497 7607 7531
rect 9321 7497 9355 7531
rect 8401 7429 8435 7463
rect 8519 7429 8553 7463
rect 5733 7361 5767 7395
rect 5917 7361 5951 7395
rect 6006 7361 6040 7395
rect 6377 7361 6411 7395
rect 7021 7361 7055 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 9505 7361 9539 7395
rect 10701 7361 10735 7395
rect 10885 7361 10919 7395
rect 11713 7361 11747 7395
rect 11989 7361 12023 7395
rect 12365 7361 12399 7395
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 8677 7293 8711 7327
rect 11529 7293 11563 7327
rect 12449 7293 12483 7327
rect 6837 7157 6871 7191
rect 10701 7157 10735 7191
rect 6285 6953 6319 6987
rect 7941 6953 7975 6987
rect 9045 6953 9079 6987
rect 9597 6953 9631 6987
rect 10517 6953 10551 6987
rect 6101 6885 6135 6919
rect 7573 6885 7607 6919
rect 9965 6885 9999 6919
rect 11345 6885 11379 6919
rect 2881 6817 2915 6851
rect 7849 6817 7883 6851
rect 10057 6817 10091 6851
rect 11529 6817 11563 6851
rect 11989 6817 12023 6851
rect 3065 6749 3099 6783
rect 4721 6749 4755 6783
rect 4977 6749 5011 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 8585 6749 8619 6783
rect 8677 6749 8711 6783
rect 8769 6749 8803 6783
rect 9321 6749 9355 6783
rect 9413 6749 9447 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 11621 6749 11655 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12173 6749 12207 6783
rect 8953 6681 8987 6715
rect 9689 6681 9723 6715
rect 9781 6681 9815 6715
rect 10149 6681 10183 6715
rect 11069 6681 11103 6715
rect 3249 6613 3283 6647
rect 10977 6613 11011 6647
rect 12357 6613 12391 6647
rect 3525 6341 3559 6375
rect 3617 6341 3651 6375
rect 8585 6341 8619 6375
rect 11529 6341 11563 6375
rect 2625 6273 2659 6307
rect 2881 6273 2915 6307
rect 3157 6273 3191 6307
rect 3433 6273 3467 6307
rect 3801 6273 3835 6307
rect 4077 6273 4111 6307
rect 4537 6273 4571 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 8033 6273 8067 6307
rect 9597 6273 9631 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 10793 6273 10827 6307
rect 11253 6273 11287 6307
rect 4261 6205 4295 6239
rect 8953 6205 8987 6239
rect 13277 6205 13311 6239
rect 2973 6137 3007 6171
rect 3249 6137 3283 6171
rect 7665 6137 7699 6171
rect 9137 6137 9171 6171
rect 9505 6137 9539 6171
rect 1501 6069 1535 6103
rect 3893 6069 3927 6103
rect 4445 6069 4479 6103
rect 7113 6069 7147 6103
rect 9045 6069 9079 6103
rect 4353 5865 4387 5899
rect 8125 5865 8159 5899
rect 8677 5865 8711 5899
rect 9781 5865 9815 5899
rect 11713 5865 11747 5899
rect 7849 5797 7883 5831
rect 12081 5797 12115 5831
rect 2237 5729 2271 5763
rect 6469 5729 6503 5763
rect 8309 5729 8343 5763
rect 9873 5729 9907 5763
rect 2145 5661 2179 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 6377 5661 6411 5695
rect 8217 5661 8251 5695
rect 8493 5661 8527 5695
rect 8953 5663 8987 5697
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9781 5661 9815 5695
rect 10333 5661 10367 5695
rect 13461 5661 13495 5695
rect 2504 5593 2538 5627
rect 3985 5593 4019 5627
rect 6714 5593 6748 5627
rect 10578 5593 10612 5627
rect 13194 5593 13228 5627
rect 1961 5525 1995 5559
rect 3617 5525 3651 5559
rect 5089 5525 5123 5559
rect 9689 5525 9723 5559
rect 10149 5525 10183 5559
rect 2973 5321 3007 5355
rect 4445 5321 4479 5355
rect 5089 5321 5123 5355
rect 7665 5321 7699 5355
rect 10425 5321 10459 5355
rect 10901 5321 10935 5355
rect 11897 5321 11931 5355
rect 13461 5321 13495 5355
rect 3433 5253 3467 5287
rect 3525 5253 3559 5287
rect 6377 5253 6411 5287
rect 7849 5253 7883 5287
rect 8953 5253 8987 5287
rect 10701 5253 10735 5287
rect 12348 5253 12382 5287
rect 1501 5185 1535 5219
rect 1768 5185 1802 5219
rect 3157 5185 3191 5219
rect 3249 5185 3283 5219
rect 3617 5185 3651 5219
rect 4629 5185 4663 5219
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 5549 5185 5583 5219
rect 5733 5185 5767 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 7021 5185 7055 5219
rect 7297 5185 7331 5219
rect 8033 5185 8067 5219
rect 8125 5185 8159 5219
rect 8493 5185 8527 5219
rect 8769 5185 8803 5219
rect 9229 5185 9263 5219
rect 9413 5185 9447 5219
rect 9873 5185 9907 5219
rect 10057 5185 10091 5219
rect 10609 5185 10643 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 5365 5117 5399 5151
rect 6837 5117 6871 5151
rect 3801 5049 3835 5083
rect 6377 5049 6411 5083
rect 11529 5049 11563 5083
rect 2881 4981 2915 5015
rect 8309 4981 8343 5015
rect 8677 4981 8711 5015
rect 9137 4981 9171 5015
rect 9413 4981 9447 5015
rect 10057 4981 10091 5015
rect 10885 4981 10919 5015
rect 11069 4981 11103 5015
rect 9781 4709 9815 4743
rect 4169 4641 4203 4675
rect 10149 4641 10183 4675
rect 3985 4573 4019 4607
rect 4997 4573 5031 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 5733 4573 5767 4607
rect 5825 4573 5859 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 9965 4573 9999 4607
rect 11161 4573 11195 4607
rect 5181 4505 5215 4539
rect 8493 4505 8527 4539
rect 9597 4505 9631 4539
rect 9781 4505 9815 4539
rect 10149 4505 10183 4539
rect 3801 4437 3835 4471
rect 5549 4437 5583 4471
rect 6009 4437 6043 4471
rect 8217 4437 8251 4471
rect 11345 4437 11379 4471
rect 3433 4233 3467 4267
rect 8401 4233 8435 4267
rect 9597 4233 9631 4267
rect 11069 4233 11103 4267
rect 3065 4165 3099 4199
rect 3709 4165 3743 4199
rect 4353 4165 4387 4199
rect 8677 4165 8711 4199
rect 2881 4097 2915 4131
rect 3157 4097 3191 4131
rect 3249 4097 3283 4131
rect 3525 4097 3559 4131
rect 3801 4097 3835 4131
rect 3893 4097 3927 4131
rect 4169 4097 4203 4131
rect 4445 4097 4479 4131
rect 4537 4097 4571 4131
rect 5069 4097 5103 4131
rect 6561 4097 6595 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 8861 4097 8895 4131
rect 9413 4097 9447 4131
rect 9689 4097 9723 4131
rect 9956 4097 9990 4131
rect 11529 4097 11563 4131
rect 11785 4097 11819 4131
rect 4813 4029 4847 4063
rect 6377 4029 6411 4063
rect 9137 4029 9171 4063
rect 6193 3961 6227 3995
rect 4077 3893 4111 3927
rect 4721 3893 4755 3927
rect 6745 3893 6779 3927
rect 8033 3893 8067 3927
rect 9045 3893 9079 3927
rect 9229 3893 9263 3927
rect 12909 3893 12943 3927
rect 4445 3689 4479 3723
rect 5549 3689 5583 3723
rect 10149 3689 10183 3723
rect 13461 3689 13495 3723
rect 3617 3621 3651 3655
rect 4169 3553 4203 3587
rect 4905 3553 4939 3587
rect 7021 3553 7055 3587
rect 7389 3553 7423 3587
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 7297 3485 7331 3519
rect 7656 3485 7690 3519
rect 10425 3485 10459 3519
rect 12081 3485 12115 3519
rect 2504 3417 2538 3451
rect 5273 3417 5307 3451
rect 6754 3417 6788 3451
rect 12348 3417 12382 3451
rect 2145 3349 2179 3383
rect 3801 3349 3835 3383
rect 5641 3349 5675 3383
rect 7113 3349 7147 3383
rect 8769 3349 8803 3383
rect 10609 3349 10643 3383
rect 3709 3145 3743 3179
rect 4813 3145 4847 3179
rect 6561 3145 6595 3179
rect 2237 3009 2271 3043
rect 2493 3009 2527 3043
rect 3893 3009 3927 3043
rect 5937 3009 5971 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 8217 3009 8251 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 8861 3009 8895 3043
rect 10066 3009 10100 3043
rect 10333 3009 10367 3043
rect 8493 2873 8527 2907
rect 8585 2873 8619 2907
rect 3617 2805 3651 2839
rect 8953 2805 8987 2839
rect 9137 2601 9171 2635
rect 9597 2601 9631 2635
rect 13461 2601 13495 2635
rect 9781 2533 9815 2567
rect 1593 2397 1627 2431
rect 2421 2397 2455 2431
rect 3617 2397 3651 2431
rect 4813 2397 4847 2431
rect 6009 2397 6043 2431
rect 7205 2397 7239 2431
rect 8401 2397 8435 2431
rect 9413 2397 9447 2431
rect 9505 2397 9539 2431
rect 9965 2397 9999 2431
rect 10793 2397 10827 2431
rect 11989 2397 12023 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 9137 2329 9171 2363
rect 9321 2329 9355 2363
rect 1409 2261 1443 2295
rect 2237 2261 2271 2295
rect 3433 2261 3467 2295
rect 4629 2261 4663 2295
rect 5825 2261 5859 2295
rect 7021 2261 7055 2295
rect 8217 2261 8251 2295
rect 10609 2261 10643 2295
rect 11805 2261 11839 2295
rect 13001 2261 13035 2295
<< metal1 >>
rect 1104 14714 13984 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13984 14714
rect 1104 14640 13984 14662
rect 934 14560 940 14612
rect 992 14600 998 14612
rect 1397 14603 1455 14609
rect 1397 14600 1409 14603
rect 992 14572 1409 14600
rect 992 14560 998 14572
rect 1397 14569 1409 14572
rect 1443 14569 1455 14603
rect 1397 14563 1455 14569
rect 2041 14603 2099 14609
rect 2041 14569 2053 14603
rect 2087 14600 2099 14603
rect 2314 14600 2320 14612
rect 2087 14572 2320 14600
rect 2087 14569 2099 14572
rect 2041 14563 2099 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 3050 14560 3056 14612
rect 3108 14560 3114 14612
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 4028 14572 4077 14600
rect 4028 14560 4034 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 5074 14560 5080 14612
rect 5132 14560 5138 14612
rect 5994 14560 6000 14612
rect 6052 14600 6058 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 6052 14572 6377 14600
rect 6052 14560 6058 14572
rect 6365 14569 6377 14572
rect 6411 14569 6423 14603
rect 6365 14563 6423 14569
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 7064 14572 7113 14600
rect 7064 14560 7070 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7101 14563 7159 14569
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7892 14572 8125 14600
rect 7892 14560 7898 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 9088 14572 9137 14600
rect 9088 14560 9094 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 3510 14492 3516 14544
rect 3568 14532 3574 14544
rect 5442 14532 5448 14544
rect 3568 14504 5448 14532
rect 3568 14492 3574 14504
rect 5442 14492 5448 14504
rect 5500 14532 5506 14544
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 5500 14504 13369 14532
rect 5500 14492 5506 14504
rect 13357 14501 13369 14504
rect 13403 14501 13415 14535
rect 13357 14495 13415 14501
rect 1578 14356 1584 14408
rect 1636 14356 1642 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2774 14396 2780 14408
rect 2271 14368 2780 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 4246 14356 4252 14408
rect 4304 14356 4310 14408
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 3694 14288 3700 14340
rect 3752 14328 3758 14340
rect 5276 14328 5304 14359
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 5408 14368 6561 14396
rect 5408 14356 5414 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7300 14328 7328 14359
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7800 14368 8309 14396
rect 7800 14356 7806 14368
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8297 14359 8355 14365
rect 8588 14368 9321 14396
rect 3752 14300 5304 14328
rect 5644 14300 7328 14328
rect 3752 14288 3758 14300
rect 5644 14272 5672 14300
rect 8588 14272 8616 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 11112 14368 11161 14396
rect 11112 14356 11118 14368
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 12124 14368 12357 14396
rect 12124 14356 12130 14368
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13136 14368 13185 14396
rect 13136 14356 13142 14368
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 5626 14220 5632 14272
rect 5684 14220 5690 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 8570 14260 8576 14272
rect 6972 14232 8576 14260
rect 6972 14220 6978 14232
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 11330 14220 11336 14272
rect 11388 14220 11394 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 11940 14232 12173 14260
rect 11940 14220 11946 14232
rect 12161 14229 12173 14232
rect 12207 14229 12219 14263
rect 12161 14223 12219 14229
rect 1104 14170 13984 14192
rect 1104 14118 4918 14170
rect 4970 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 5238 14170
rect 5290 14118 10918 14170
rect 10970 14118 10982 14170
rect 11034 14118 11046 14170
rect 11098 14118 11110 14170
rect 11162 14118 11174 14170
rect 11226 14118 11238 14170
rect 11290 14118 13984 14170
rect 1104 14096 13984 14118
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 2884 14028 3525 14056
rect 2884 13932 2912 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 4525 14059 4583 14065
rect 4525 14056 4537 14059
rect 3513 14019 3571 14025
rect 4172 14028 4537 14056
rect 4172 13997 4200 14028
rect 4525 14025 4537 14028
rect 4571 14025 4583 14059
rect 4525 14019 4583 14025
rect 6914 14016 6920 14068
rect 6972 14016 6978 14068
rect 3605 13991 3663 13997
rect 3605 13988 3617 13991
rect 2976 13960 3617 13988
rect 2976 13932 3004 13960
rect 3605 13957 3617 13960
rect 3651 13988 3663 13991
rect 4157 13991 4215 13997
rect 4157 13988 4169 13991
rect 3651 13960 4169 13988
rect 3651 13957 3663 13960
rect 3605 13951 3663 13957
rect 4157 13957 4169 13960
rect 4203 13957 4215 13991
rect 4430 13988 4436 14000
rect 4157 13951 4215 13957
rect 4264 13960 4436 13988
rect 2866 13880 2872 13932
rect 2924 13880 2930 13932
rect 2958 13880 2964 13932
rect 3016 13880 3022 13932
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 3510 13920 3516 13932
rect 3283 13892 3516 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 3712 13852 3740 13883
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3844 13892 3985 13920
rect 3844 13880 3850 13892
rect 3973 13889 3985 13892
rect 4019 13920 4031 13923
rect 4062 13920 4068 13932
rect 4019 13892 4068 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4264 13929 4292 13960
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 5350 13988 5356 14000
rect 4540 13960 5356 13988
rect 4540 13932 4568 13960
rect 5350 13948 5356 13960
rect 5408 13948 5414 14000
rect 6932 13963 6960 14016
rect 6917 13957 6975 13963
rect 6644 13945 6702 13951
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4522 13920 4528 13932
rect 4387 13892 4528 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4663 13892 4844 13920
rect 6644 13911 6656 13945
rect 6690 13911 6702 13945
rect 6644 13905 6702 13911
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4816 13852 4844 13892
rect 6656 13864 6684 13905
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 6917 13923 6929 13957
rect 6963 13923 6975 13957
rect 7098 13948 7104 14000
rect 7156 13948 7162 14000
rect 7285 13991 7343 13997
rect 7285 13957 7297 13991
rect 7331 13988 7343 13991
rect 7742 13988 7748 14000
rect 7331 13960 7748 13988
rect 7331 13957 7343 13960
rect 7285 13951 7343 13957
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 9048 13960 10180 13988
rect 6917 13917 6975 13923
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13910 7067 13923
rect 7190 13920 7196 13932
rect 7116 13910 7196 13920
rect 7055 13892 7196 13910
rect 7055 13889 7144 13892
rect 7009 13883 7144 13889
rect 7024 13882 7144 13883
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 8662 13880 8668 13932
rect 8720 13920 8726 13932
rect 9048 13929 9076 13960
rect 10152 13932 10180 13960
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8720 13892 9045 13920
rect 8720 13880 8726 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9033 13883 9091 13889
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9766 13920 9772 13932
rect 9263 13892 9772 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 10192 13892 10701 13920
rect 10192 13880 10198 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10870 13880 10876 13932
rect 10928 13880 10934 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11514 13920 11520 13932
rect 11011 13892 11520 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 3712 13824 4844 13852
rect 4816 13796 4844 13824
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 9125 13855 9183 13861
rect 6880 13824 6960 13852
rect 6880 13812 6886 13824
rect 4341 13787 4399 13793
rect 4341 13784 4353 13787
rect 3344 13756 4353 13784
rect 3234 13676 3240 13728
rect 3292 13676 3298 13728
rect 3344 13725 3372 13756
rect 4341 13753 4353 13756
rect 4387 13753 4399 13787
rect 4341 13747 4399 13753
rect 4798 13744 4804 13796
rect 4856 13744 4862 13796
rect 6932 13793 6960 13824
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9674 13852 9680 13864
rect 9171 13824 9680 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 6917 13787 6975 13793
rect 6917 13753 6929 13787
rect 6963 13753 6975 13787
rect 6917 13747 6975 13753
rect 3329 13719 3387 13725
rect 3329 13685 3341 13719
rect 3375 13685 3387 13719
rect 3329 13679 3387 13685
rect 3970 13676 3976 13728
rect 4028 13676 4034 13728
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 6236 13688 7297 13716
rect 6236 13676 6242 13688
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 10686 13676 10692 13728
rect 10744 13676 10750 13728
rect 1104 13626 13984 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13984 13626
rect 1104 13552 13984 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 3970 13512 3976 13524
rect 3467 13484 3976 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4120 13484 5181 13512
rect 4120 13472 4126 13484
rect 5169 13481 5181 13484
rect 5215 13512 5227 13515
rect 5626 13512 5632 13524
rect 5215 13484 5632 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6178 13472 6184 13524
rect 6236 13472 6242 13524
rect 6270 13472 6276 13524
rect 6328 13472 6334 13524
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6730 13512 6736 13524
rect 6420 13484 6736 13512
rect 6420 13472 6426 13484
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 6822 13472 6828 13524
rect 6880 13472 6886 13524
rect 8662 13512 8668 13524
rect 6932 13484 8668 13512
rect 2869 13447 2927 13453
rect 2869 13413 2881 13447
rect 2915 13444 2927 13447
rect 3050 13444 3056 13456
rect 2915 13416 3056 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3050 13404 3056 13416
rect 3108 13444 3114 13456
rect 3694 13444 3700 13456
rect 3108 13416 3700 13444
rect 3108 13404 3114 13416
rect 3694 13404 3700 13416
rect 3752 13404 3758 13456
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 5537 13447 5595 13453
rect 5537 13444 5549 13447
rect 5500 13416 5549 13444
rect 5500 13404 5506 13416
rect 5537 13413 5549 13416
rect 5583 13444 5595 13447
rect 6932 13444 6960 13484
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 5583 13416 6960 13444
rect 5583 13413 5595 13416
rect 5537 13407 5595 13413
rect 3789 13379 3847 13385
rect 3789 13376 3801 13379
rect 2700 13348 3801 13376
rect 2700 13320 2728 13348
rect 3789 13345 3801 13348
rect 3835 13345 3847 13379
rect 3789 13339 3847 13345
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13308 1547 13311
rect 2682 13308 2688 13320
rect 1535 13280 2688 13308
rect 1535 13277 1547 13280
rect 1489 13271 1547 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3326 13308 3332 13320
rect 3099 13280 3332 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13300 3571 13311
rect 5460 13308 5488 13404
rect 6178 13336 6184 13388
rect 6236 13336 6242 13388
rect 3620 13300 5488 13308
rect 3559 13280 5488 13300
rect 3559 13277 3648 13280
rect 3513 13272 3648 13277
rect 3513 13271 3571 13272
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5776 13280 5825 13308
rect 5776 13268 5782 13280
rect 5813 13277 5825 13280
rect 5859 13308 5871 13311
rect 6196 13308 6224 13336
rect 6288 13317 6316 13416
rect 6730 13376 6736 13388
rect 6472 13348 6736 13376
rect 6472 13317 6500 13348
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 6932 13317 6960 13416
rect 5859 13280 6224 13308
rect 6273 13311 6331 13317
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 10054 13311 10112 13317
rect 10054 13308 10066 13311
rect 9732 13280 10066 13308
rect 9732 13268 9738 13280
rect 10054 13277 10066 13280
rect 10100 13277 10112 13311
rect 10054 13271 10112 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10367 13280 10425 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10413 13277 10425 13280
rect 10459 13308 10471 13311
rect 12066 13308 12072 13320
rect 10459 13280 12072 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 1756 13243 1814 13249
rect 1756 13209 1768 13243
rect 1802 13240 1814 13243
rect 2130 13240 2136 13252
rect 1802 13212 2136 13240
rect 1802 13209 1814 13212
rect 1756 13203 1814 13209
rect 2130 13200 2136 13212
rect 2188 13200 2194 13252
rect 4034 13243 4092 13249
rect 4034 13240 4046 13243
rect 2884 13212 3280 13240
rect 2884 13184 2912 13212
rect 2866 13132 2872 13184
rect 2924 13132 2930 13184
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 3252 13181 3280 13212
rect 3804 13212 4046 13240
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 3016 13144 3157 13172
rect 3016 13132 3022 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13141 3295 13175
rect 3237 13135 3295 13141
rect 3513 13175 3571 13181
rect 3513 13141 3525 13175
rect 3559 13172 3571 13175
rect 3804 13172 3832 13212
rect 4034 13209 4046 13212
rect 4080 13209 4092 13243
rect 4034 13203 4092 13209
rect 5350 13200 5356 13252
rect 5408 13200 5414 13252
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 6362 13240 6368 13252
rect 5951 13212 6368 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 6362 13200 6368 13212
rect 6420 13240 6426 13252
rect 10686 13249 10692 13252
rect 6549 13243 6607 13249
rect 6549 13240 6561 13243
rect 6420 13212 6561 13240
rect 6420 13200 6426 13212
rect 6549 13209 6561 13212
rect 6595 13209 6607 13243
rect 7438 13243 7496 13249
rect 7438 13240 7450 13243
rect 6549 13203 6607 13209
rect 6932 13212 7450 13240
rect 3559 13144 3832 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 3936 13144 6009 13172
rect 3936 13132 3942 13144
rect 5997 13141 6009 13144
rect 6043 13172 6055 13175
rect 6454 13172 6460 13184
rect 6043 13144 6460 13172
rect 6043 13141 6055 13144
rect 5997 13135 6055 13141
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 6932 13181 6960 13212
rect 7438 13209 7450 13212
rect 7484 13209 7496 13243
rect 10680 13240 10692 13249
rect 10647 13212 10692 13240
rect 7438 13203 7496 13209
rect 10680 13203 10692 13212
rect 10686 13200 10692 13203
rect 10744 13200 10750 13252
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13141 6975 13175
rect 6917 13135 6975 13141
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 11790 13172 11796 13184
rect 9272 13144 11796 13172
rect 9272 13132 9278 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 1104 13082 13984 13104
rect 1104 13030 4918 13082
rect 4970 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 5238 13082
rect 5290 13030 10918 13082
rect 10970 13030 10982 13082
rect 11034 13030 11046 13082
rect 11098 13030 11110 13082
rect 11162 13030 11174 13082
rect 11226 13030 11238 13082
rect 11290 13030 13984 13082
rect 1104 13008 13984 13030
rect 2130 12928 2136 12980
rect 2188 12928 2194 12980
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 3878 12968 3884 12980
rect 2924 12940 3884 12968
rect 2924 12928 2930 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4580 12940 4629 12968
rect 4580 12928 4586 12940
rect 4617 12937 4629 12940
rect 4663 12937 4675 12971
rect 4617 12931 4675 12937
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 4893 12971 4951 12977
rect 4893 12968 4905 12971
rect 4856 12940 4905 12968
rect 4856 12928 4862 12940
rect 4893 12937 4905 12940
rect 4939 12937 4951 12971
rect 5810 12968 5816 12980
rect 4893 12931 4951 12937
rect 5184 12940 5816 12968
rect 5061 12903 5119 12909
rect 3252 12872 3648 12900
rect 2314 12792 2320 12844
rect 2372 12792 2378 12844
rect 3252 12841 3280 12872
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 2746 12804 3249 12832
rect 2746 12776 2774 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3493 12835 3551 12841
rect 3493 12832 3505 12835
rect 3384 12804 3505 12832
rect 3384 12792 3390 12804
rect 3493 12801 3505 12804
rect 3539 12801 3551 12835
rect 3620 12832 3648 12872
rect 5061 12869 5073 12903
rect 5107 12900 5119 12903
rect 5184 12900 5212 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7800 12940 7941 12968
rect 7800 12928 7806 12940
rect 7929 12937 7941 12940
rect 7975 12937 7987 12971
rect 7929 12931 7987 12937
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 9766 12968 9772 12980
rect 9723 12940 9772 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 9858 12928 9864 12980
rect 9916 12928 9922 12980
rect 11514 12928 11520 12980
rect 11572 12928 11578 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11848 12940 12173 12968
rect 11848 12928 11854 12940
rect 12161 12937 12173 12940
rect 12207 12968 12219 12971
rect 12207 12940 12480 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 5107 12872 5212 12900
rect 5107 12869 5119 12872
rect 5061 12863 5119 12869
rect 5258 12860 5264 12912
rect 5316 12860 5322 12912
rect 7208 12900 7236 12928
rect 6564 12872 7236 12900
rect 6564 12841 6592 12872
rect 8938 12860 8944 12912
rect 8996 12860 9002 12912
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 12253 12903 12311 12909
rect 12253 12900 12265 12903
rect 10652 12872 12265 12900
rect 10652 12860 10658 12872
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 3620 12804 6561 12832
rect 3493 12795 3551 12801
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6805 12835 6863 12841
rect 6805 12832 6817 12835
rect 6549 12795 6607 12801
rect 6656 12804 6817 12832
rect 2682 12724 2688 12776
rect 2740 12736 2774 12776
rect 2740 12724 2746 12736
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6656 12764 6684 12804
rect 6805 12801 6817 12804
rect 6851 12801 6863 12835
rect 8956 12832 8984 12860
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 8956 12804 9321 12832
rect 6805 12795 6863 12801
rect 9309 12801 9321 12804
rect 9355 12832 9367 12835
rect 9490 12832 9496 12844
rect 9355 12804 9496 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9490 12792 9496 12804
rect 9548 12832 9554 12844
rect 10888 12841 10916 12872
rect 12253 12869 12265 12872
rect 12299 12869 12311 12903
rect 12452 12900 12480 12940
rect 12452 12872 12572 12900
rect 12253 12863 12311 12869
rect 9858 12835 9916 12841
rect 9858 12832 9870 12835
rect 9548 12804 9870 12832
rect 9548 12792 9554 12804
rect 9858 12801 9870 12804
rect 9904 12832 9916 12835
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 9904 12804 10701 12832
rect 9904 12801 9916 12804
rect 9858 12795 9916 12801
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11606 12832 11612 12844
rect 11195 12804 11612 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 6328 12736 6684 12764
rect 6328 12724 6334 12736
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9214 12764 9220 12776
rect 8720 12736 9220 12764
rect 8720 12724 8726 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 9784 12736 10333 12764
rect 5258 12696 5264 12708
rect 5000 12668 5264 12696
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 5000 12628 5028 12668
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 9784 12640 9812 12736
rect 10321 12733 10333 12736
rect 10367 12764 10379 12767
rect 10410 12764 10416 12776
rect 10367 12736 10416 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10980 12764 11008 12795
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 12544 12841 12572 12872
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 11701 12767 11759 12773
rect 10980 12736 11376 12764
rect 11348 12708 11376 12736
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 10781 12699 10839 12705
rect 10781 12665 10793 12699
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 4028 12600 5028 12628
rect 5077 12631 5135 12637
rect 4028 12588 4034 12600
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5350 12628 5356 12640
rect 5123 12600 5356 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 8938 12588 8944 12640
rect 8996 12588 9002 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9766 12588 9772 12640
rect 9824 12588 9830 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10275 12600 10517 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10796 12628 10824 12659
rect 11330 12656 11336 12708
rect 11388 12656 11394 12708
rect 11716 12696 11744 12727
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 12391 12736 12572 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 12544 12708 12572 12736
rect 12434 12696 12440 12708
rect 11716 12668 12440 12696
rect 12434 12656 12440 12668
rect 12492 12656 12498 12708
rect 12526 12656 12532 12708
rect 12584 12656 12590 12708
rect 12342 12628 12348 12640
rect 10796 12600 12348 12628
rect 10505 12591 10563 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12710 12588 12716 12640
rect 12768 12588 12774 12640
rect 1104 12538 13984 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13984 12538
rect 1104 12464 13984 12486
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 4632 12396 4813 12424
rect 2225 12359 2283 12365
rect 2225 12325 2237 12359
rect 2271 12356 2283 12359
rect 3694 12356 3700 12368
rect 2271 12328 3700 12356
rect 2271 12325 2283 12328
rect 2225 12319 2283 12325
rect 3694 12316 3700 12328
rect 3752 12316 3758 12368
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 4632 12288 4660 12396
rect 4801 12393 4813 12396
rect 4847 12393 4859 12427
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 4801 12387 4859 12393
rect 4908 12396 5549 12424
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 4908 12356 4936 12396
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 5537 12387 5595 12393
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 5810 12384 5816 12436
rect 5868 12384 5874 12436
rect 5994 12433 6000 12436
rect 5975 12427 6000 12433
rect 5975 12393 5987 12427
rect 5975 12387 6000 12393
rect 5994 12384 6000 12387
rect 6052 12384 6058 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6144 12396 6561 12424
rect 6144 12384 6150 12396
rect 6549 12393 6561 12396
rect 6595 12393 6607 12427
rect 6549 12387 6607 12393
rect 6730 12384 6736 12436
rect 6788 12384 6794 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 9858 12424 9864 12436
rect 9815 12396 9864 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10008 12396 11284 12424
rect 10008 12384 10014 12396
rect 11256 12368 11284 12396
rect 4764 12328 4936 12356
rect 4764 12316 4770 12328
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 9033 12359 9091 12365
rect 9033 12356 9045 12359
rect 8720 12328 9045 12356
rect 8720 12316 8726 12328
rect 9033 12325 9045 12328
rect 9079 12325 9091 12359
rect 9033 12319 9091 12325
rect 9232 12328 11100 12356
rect 4798 12288 4804 12300
rect 3016 12260 3280 12288
rect 4632 12260 4804 12288
rect 3016 12248 3022 12260
rect 3252 12232 3280 12260
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4908 12260 5856 12288
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 2498 12112 2504 12164
rect 2556 12112 2562 12164
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 2041 12087 2099 12093
rect 2041 12084 2053 12087
rect 1728 12056 2053 12084
rect 1728 12044 1734 12056
rect 2041 12053 2053 12056
rect 2087 12053 2099 12087
rect 2041 12047 2099 12053
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2648 12056 2697 12084
rect 2648 12044 2654 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2884 12084 2912 12183
rect 3068 12152 3096 12183
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 4908 12220 4936 12260
rect 5828 12232 5856 12260
rect 9232 12232 9260 12328
rect 10962 12288 10968 12300
rect 9692 12260 10272 12288
rect 9692 12232 9720 12260
rect 4800 12195 4936 12220
rect 4755 12192 4936 12195
rect 5169 12223 5227 12229
rect 4755 12189 4828 12192
rect 4246 12152 4252 12164
rect 3068 12124 4252 12152
rect 4246 12112 4252 12124
rect 4304 12152 4310 12164
rect 4755 12155 4767 12189
rect 4801 12158 4828 12189
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 5534 12220 5540 12232
rect 5215 12192 5540 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 5810 12180 5816 12232
rect 5868 12180 5874 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 5960 12192 6408 12220
rect 5960 12180 5966 12192
rect 4801 12155 4813 12158
rect 4304 12124 4660 12152
rect 4755 12149 4813 12155
rect 4985 12155 5043 12161
rect 4304 12112 4310 12124
rect 4632 12096 4660 12124
rect 4985 12121 4997 12155
rect 5031 12152 5043 12155
rect 5920 12152 5948 12180
rect 5031 12124 5948 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 6380 12161 6408 12192
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9674 12180 9680 12232
rect 9732 12180 9738 12232
rect 9950 12229 9956 12232
rect 9948 12220 9956 12229
rect 9911 12192 9956 12220
rect 9948 12183 9956 12192
rect 9950 12180 9956 12183
rect 10008 12180 10014 12232
rect 10244 12229 10272 12260
rect 10796 12260 10968 12288
rect 10244 12223 10323 12229
rect 10244 12192 10277 12223
rect 10265 12189 10277 12192
rect 10311 12189 10323 12223
rect 10265 12183 10323 12189
rect 10410 12180 10416 12232
rect 10468 12180 10474 12232
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 10796 12229 10824 12260
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 6365 12155 6423 12161
rect 6365 12121 6377 12155
rect 6411 12152 6423 12155
rect 7098 12152 7104 12164
rect 6411 12124 7104 12152
rect 6411 12121 6423 12124
rect 6365 12115 6423 12121
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 9858 12152 9864 12164
rect 9232 12124 9864 12152
rect 3050 12084 3056 12096
rect 2884 12056 3056 12084
rect 2685 12047 2743 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3510 12084 3516 12096
rect 3384 12056 3516 12084
rect 3384 12044 3390 12056
rect 3510 12044 3516 12056
rect 3568 12044 3574 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5408 12056 5549 12084
rect 5408 12044 5414 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 5971 12087 6029 12093
rect 5971 12084 5983 12087
rect 5776 12056 5983 12084
rect 5776 12044 5782 12056
rect 5971 12053 5983 12056
rect 6017 12053 6029 12087
rect 5971 12047 6029 12053
rect 6575 12087 6633 12093
rect 6575 12053 6587 12087
rect 6621 12084 6633 12087
rect 9232 12084 9260 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10042 12112 10048 12164
rect 10100 12112 10106 12164
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10594 12152 10600 12164
rect 10183 12124 10600 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 11072 12152 11100 12328
rect 11238 12316 11244 12368
rect 11296 12316 11302 12368
rect 11790 12356 11796 12368
rect 11532 12328 11796 12356
rect 11532 12297 11560 12328
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11195 12260 11529 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11756 12260 12020 12288
rect 11756 12248 11762 12260
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12220 11299 12223
rect 11330 12220 11336 12232
rect 11287 12192 11336 12220
rect 11287 12189 11299 12192
rect 11241 12183 11299 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12189 11851 12223
rect 11992 12218 12020 12260
rect 12066 12218 12072 12232
rect 11992 12190 12072 12218
rect 11793 12183 11851 12189
rect 11808 12152 11836 12183
rect 12066 12180 12072 12190
rect 12124 12180 12130 12232
rect 12336 12223 12394 12229
rect 12336 12189 12348 12223
rect 12382 12189 12394 12223
rect 12336 12183 12394 12189
rect 11072 12124 12204 12152
rect 6621 12056 9260 12084
rect 6621 12053 6633 12056
rect 6575 12047 6633 12053
rect 9306 12044 9312 12096
rect 9364 12044 9370 12096
rect 9398 12044 9404 12096
rect 9456 12044 9462 12096
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 11790 12084 11796 12096
rect 11296 12056 11796 12084
rect 11296 12044 11302 12056
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 11974 12044 11980 12096
rect 12032 12044 12038 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12176 12084 12204 12124
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 12360 12152 12388 12183
rect 12308 12124 12388 12152
rect 12308 12112 12314 12124
rect 12618 12084 12624 12096
rect 12124 12056 12624 12084
rect 12124 12044 12130 12056
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 12676 12056 13461 12084
rect 12676 12044 12682 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 1104 11994 13984 12016
rect 1104 11942 4918 11994
rect 4970 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 5238 11994
rect 5290 11942 10918 11994
rect 10970 11942 10982 11994
rect 11034 11942 11046 11994
rect 11098 11942 11110 11994
rect 11162 11942 11174 11994
rect 11226 11942 11238 11994
rect 11290 11942 13984 11994
rect 1104 11920 13984 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 2556 11852 2973 11880
rect 2556 11840 2562 11852
rect 2961 11849 2973 11852
rect 3007 11849 3019 11883
rect 2961 11843 3019 11849
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3467 11852 3501 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 2682 11812 2688 11824
rect 1504 11784 2688 11812
rect 1504 11753 1532 11784
rect 2682 11772 2688 11784
rect 2740 11772 2746 11824
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 3436 11812 3464 11843
rect 3694 11840 3700 11892
rect 3752 11840 3758 11892
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4488 11852 4813 11880
rect 4488 11840 4494 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11849 5135 11883
rect 5077 11843 5135 11849
rect 4709 11815 4767 11821
rect 3292 11784 4108 11812
rect 3292 11772 3298 11784
rect 1762 11753 1768 11756
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 1756 11707 1768 11753
rect 1762 11704 1768 11707
rect 1820 11704 1826 11756
rect 4080 11753 4108 11784
rect 4479 11781 4537 11787
rect 4479 11756 4491 11781
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3513 11747 3571 11753
rect 3191 11716 3372 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3344 11688 3372 11716
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 4065 11747 4123 11753
rect 3559 11716 4016 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 2924 11648 3249 11676
rect 2924 11636 2930 11648
rect 3237 11645 3249 11648
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 3326 11636 3332 11688
rect 3384 11636 3390 11688
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3988 11685 4016 11716
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4430 11704 4436 11756
rect 4488 11747 4491 11756
rect 4525 11778 4537 11781
rect 4709 11781 4721 11815
rect 4755 11812 4767 11815
rect 4890 11812 4896 11824
rect 4755 11784 4896 11812
rect 4755 11781 4767 11784
rect 4525 11747 4552 11778
rect 4709 11775 4767 11781
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 4982 11772 4988 11824
rect 5040 11772 5046 11824
rect 5092 11812 5120 11843
rect 5166 11840 5172 11892
rect 5224 11840 5230 11892
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5408 11852 6377 11880
rect 5408 11840 5414 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6365 11843 6423 11849
rect 6748 11852 7021 11880
rect 5721 11815 5779 11821
rect 5092 11784 5212 11812
rect 4488 11716 4552 11747
rect 4488 11704 4494 11716
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 3660 11648 3893 11676
rect 3660 11636 3666 11648
rect 3881 11645 3893 11648
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4246 11676 4252 11688
rect 4203 11648 4252 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 3988 11608 4016 11639
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 4798 11636 4804 11688
rect 4856 11636 4862 11688
rect 4908 11676 4936 11772
rect 5074 11676 5080 11688
rect 4908 11648 5080 11676
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 5184 11676 5212 11784
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 5994 11812 6000 11824
rect 5767 11784 6000 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 6748 11821 6776 11852
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 7009 11843 7067 11849
rect 8036 11852 8493 11880
rect 8036 11821 8064 11852
rect 8481 11849 8493 11852
rect 8527 11849 8539 11883
rect 8481 11843 8539 11849
rect 10318 11840 10324 11892
rect 10376 11840 10382 11892
rect 10413 11883 10471 11889
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 10686 11880 10692 11892
rect 10459 11852 10692 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 10686 11840 10692 11852
rect 10744 11840 10750 11892
rect 10778 11840 10784 11892
rect 10836 11840 10842 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10928 11852 11161 11880
rect 10928 11840 10934 11852
rect 11149 11849 11161 11852
rect 11195 11880 11207 11883
rect 11330 11880 11336 11892
rect 11195 11852 11336 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11606 11840 11612 11892
rect 11664 11840 11670 11892
rect 11790 11840 11796 11892
rect 11848 11840 11854 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12216 11852 12388 11880
rect 12216 11840 12222 11852
rect 6517 11815 6575 11821
rect 6517 11781 6529 11815
rect 6563 11812 6575 11815
rect 6733 11815 6791 11821
rect 6563 11781 6592 11812
rect 6517 11775 6592 11781
rect 6733 11781 6745 11815
rect 6779 11781 6791 11815
rect 7469 11815 7527 11821
rect 7469 11812 7481 11815
rect 6733 11775 6791 11781
rect 6840 11784 7481 11812
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 5859 11716 6500 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 5445 11679 5503 11685
rect 5445 11676 5457 11679
rect 5184 11648 5457 11676
rect 5445 11645 5457 11648
rect 5491 11676 5503 11679
rect 6086 11676 6092 11688
rect 5491 11648 6092 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 4341 11611 4399 11617
rect 4341 11608 4353 11611
rect 3988 11580 4353 11608
rect 4341 11577 4353 11580
rect 4387 11608 4399 11611
rect 4724 11608 4752 11636
rect 4387 11580 4752 11608
rect 4816 11608 4844 11636
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 4816 11580 5365 11608
rect 4387 11577 4399 11580
rect 4341 11571 4399 11577
rect 5353 11577 5365 11580
rect 5399 11577 5411 11611
rect 5353 11571 5411 11577
rect 5997 11611 6055 11617
rect 5997 11577 6009 11611
rect 6043 11608 6055 11611
rect 6270 11608 6276 11620
rect 6043 11580 6276 11608
rect 6043 11577 6055 11580
rect 5997 11571 6055 11577
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2869 11543 2927 11549
rect 2869 11540 2881 11543
rect 2832 11512 2881 11540
rect 2832 11500 2838 11512
rect 2869 11509 2881 11512
rect 2915 11540 2927 11543
rect 4246 11540 4252 11552
rect 2915 11512 4252 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 5810 11540 5816 11552
rect 4571 11512 5816 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 5810 11500 5816 11512
rect 5868 11540 5874 11552
rect 6012 11540 6040 11571
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 6472 11552 6500 11716
rect 6564 11688 6592 11775
rect 6840 11688 6868 11784
rect 7469 11781 7481 11784
rect 7515 11781 7527 11815
rect 7469 11775 7527 11781
rect 8021 11815 8079 11821
rect 8021 11781 8033 11815
rect 8067 11781 8079 11815
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 8021 11775 8079 11781
rect 8128 11784 9137 11812
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 8128 11744 8156 11784
rect 9125 11781 9137 11784
rect 9171 11812 9183 11815
rect 9398 11812 9404 11824
rect 9171 11784 9404 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9398 11772 9404 11784
rect 9456 11772 9462 11824
rect 9766 11812 9772 11824
rect 9508 11784 9772 11812
rect 7239 11716 8156 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7484 11688 7512 11716
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 9508 11753 9536 11784
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 10229 11815 10287 11821
rect 10229 11781 10241 11815
rect 10275 11812 10287 11815
rect 10336 11812 10364 11840
rect 11808 11812 11836 11840
rect 10275 11784 11560 11812
rect 10275 11781 10287 11784
rect 10229 11775 10287 11781
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9640 11716 9689 11744
rect 9640 11704 9646 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10137 11747 10195 11753
rect 10137 11744 10149 11747
rect 10100 11716 10149 11744
rect 10100 11704 10106 11716
rect 10137 11713 10149 11716
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11744 10747 11747
rect 10735 11716 10916 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 6822 11636 6828 11688
rect 6880 11636 6886 11688
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9306 11676 9312 11688
rect 8895 11648 9312 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9306 11636 9312 11648
rect 9364 11676 9370 11688
rect 10336 11676 10364 11704
rect 9364 11648 10364 11676
rect 10413 11679 10471 11685
rect 9364 11636 9370 11648
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7834 11608 7840 11620
rect 6972 11580 7840 11608
rect 6972 11568 6978 11580
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 10428 11608 10456 11639
rect 9968 11580 10456 11608
rect 10888 11608 10916 11716
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 11238 11704 11244 11756
rect 11296 11704 11302 11756
rect 11532 11753 11560 11784
rect 11716 11784 11836 11812
rect 11716 11753 11744 11784
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11992 11744 12020 11840
rect 12250 11772 12256 11824
rect 12308 11772 12314 11824
rect 12360 11821 12388 11852
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12492 11852 12725 11880
rect 12492 11840 12498 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 12345 11815 12403 11821
rect 12345 11781 12357 11815
rect 12391 11781 12403 11815
rect 12345 11775 12403 11781
rect 12618 11772 12624 11824
rect 12676 11812 12682 11824
rect 12676 11784 13032 11812
rect 12676 11772 12682 11784
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11992 11716 12081 11744
rect 11885 11707 11943 11713
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 10980 11676 11008 11704
rect 11808 11676 11836 11707
rect 10980 11648 11836 11676
rect 11238 11608 11244 11620
rect 10888 11580 11244 11608
rect 9968 11552 9996 11580
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 11606 11608 11612 11620
rect 11388 11580 11612 11608
rect 11388 11568 11394 11580
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 11900 11608 11928 11707
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 13004 11753 13032 11784
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 12544 11676 12572 11707
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12544 11648 12909 11676
rect 12544 11608 12572 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 11900 11580 12572 11608
rect 5868 11512 6040 11540
rect 5868 11500 5874 11512
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6512 11512 6561 11540
rect 6512 11500 6518 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6549 11503 6607 11509
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7064 11512 7389 11540
rect 7064 11500 7070 11512
rect 7377 11509 7389 11512
rect 7423 11540 7435 11543
rect 8662 11540 8668 11552
rect 7423 11512 8668 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9214 11540 9220 11552
rect 9079 11512 9220 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9950 11540 9956 11552
rect 9732 11512 9956 11540
rect 9732 11500 9738 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10962 11540 10968 11552
rect 10468 11512 10968 11540
rect 10468 11500 10474 11512
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 12158 11540 12164 11552
rect 11112 11512 12164 11540
rect 11112 11500 11118 11512
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 1104 11450 13984 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13984 11450
rect 1104 11376 13984 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2372 11308 2421 11336
rect 2372 11296 2378 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 2590 11296 2596 11348
rect 2648 11296 2654 11348
rect 4338 11336 4344 11348
rect 3896 11308 4344 11336
rect 2225 11271 2283 11277
rect 2225 11237 2237 11271
rect 2271 11268 2283 11271
rect 2608 11268 2636 11296
rect 3326 11268 3332 11280
rect 2271 11240 2636 11268
rect 2700 11240 3332 11268
rect 2271 11237 2283 11240
rect 2225 11231 2283 11237
rect 1670 11160 1676 11212
rect 1728 11160 1734 11212
rect 2700 11209 2728 11240
rect 3326 11228 3332 11240
rect 3384 11228 3390 11280
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 3108 11172 3157 11200
rect 3108 11160 3114 11172
rect 3145 11169 3157 11172
rect 3191 11200 3203 11203
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 3191 11172 3801 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3789 11163 3847 11169
rect 1688 11132 1716 11160
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1688 11104 1869 11132
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 2915 11135 2973 11141
rect 2915 11101 2927 11135
rect 2961 11132 2973 11135
rect 3896 11132 3924 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 5166 11336 5172 11348
rect 4479 11308 5172 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4890 11268 4896 11280
rect 4028 11240 4896 11268
rect 4028 11228 4034 11240
rect 4890 11228 4896 11240
rect 4948 11228 4954 11280
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4571 11172 4936 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4908 11144 4936 11172
rect 2961 11104 3924 11132
rect 4065 11135 4123 11141
rect 2961 11101 2973 11104
rect 2915 11095 2973 11101
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4338 11132 4344 11144
rect 4111 11104 4344 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2501 11067 2559 11073
rect 2501 11064 2513 11067
rect 1995 11036 2513 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 2501 11033 2513 11036
rect 2547 11033 2559 11067
rect 2501 11027 2559 11033
rect 2792 10996 2820 11095
rect 4338 11092 4344 11104
rect 4396 11132 4402 11144
rect 4706 11132 4712 11144
rect 4396 11104 4712 11132
rect 4396 11092 4402 11104
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 5000 11141 5028 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6362 11336 6368 11348
rect 6319 11308 6368 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6546 11296 6552 11348
rect 6604 11296 6610 11348
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 7098 11296 7104 11348
rect 7156 11296 7162 11348
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7742 11336 7748 11348
rect 7423 11308 7748 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7742 11296 7748 11308
rect 7800 11336 7806 11348
rect 8389 11339 8447 11345
rect 8389 11336 8401 11339
rect 7800 11308 8401 11336
rect 7800 11296 7806 11308
rect 8389 11305 8401 11308
rect 8435 11336 8447 11339
rect 8938 11336 8944 11348
rect 8435 11308 8944 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 5626 11268 5632 11280
rect 5092 11240 5632 11268
rect 5092 11144 5120 11240
rect 5626 11228 5632 11240
rect 5684 11268 5690 11280
rect 6564 11268 6592 11296
rect 5684 11240 6592 11268
rect 5684 11228 5690 11240
rect 5902 11200 5908 11212
rect 5276 11172 5908 11200
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 3053 11067 3111 11073
rect 3053 11033 3065 11067
rect 3099 11064 3111 11067
rect 3234 11064 3240 11076
rect 3099 11036 3240 11064
rect 3099 11033 3111 11036
rect 3053 11027 3111 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 4617 11067 4675 11073
rect 4617 11064 4629 11067
rect 4080 11036 4629 11064
rect 4080 11008 4108 11036
rect 4617 11033 4629 11036
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 2866 10996 2872 11008
rect 2792 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 4062 10956 4068 11008
rect 4120 10956 4126 11008
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4706 10996 4712 11008
rect 4295 10968 4712 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 5000 10996 5028 11095
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5276 11141 5304 11172
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6178 11200 6184 11212
rect 6052 11172 6184 11200
rect 6052 11160 6058 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 5626 11092 5632 11144
rect 5684 11092 5690 11144
rect 6380 11141 6408 11240
rect 6932 11200 6960 11296
rect 7466 11228 7472 11280
rect 7524 11228 7530 11280
rect 7650 11228 7656 11280
rect 7708 11268 7714 11280
rect 7929 11271 7987 11277
rect 7929 11268 7941 11271
rect 7708 11240 7941 11268
rect 7708 11228 7714 11240
rect 7929 11237 7941 11240
rect 7975 11237 7987 11271
rect 7929 11231 7987 11237
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 6840 11172 6960 11200
rect 7760 11172 8217 11200
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6730 11132 6736 11144
rect 6687 11104 6736 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6840 11141 6868 11172
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 6963 11104 7573 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7300 11076 7328 11104
rect 7561 11101 7573 11104
rect 7607 11132 7619 11135
rect 7760 11132 7788 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 7607 11104 7788 11132
rect 7837 11135 7895 11141
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 7926 11132 7932 11144
rect 7883 11104 7932 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8294 11132 8300 11144
rect 8159 11104 8300 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8496 11141 8524 11308
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10652 11308 11376 11336
rect 10652 11296 10658 11308
rect 8662 11228 8668 11280
rect 8720 11228 8726 11280
rect 11238 11228 11244 11280
rect 11296 11228 11302 11280
rect 11348 11268 11376 11308
rect 11422 11296 11428 11348
rect 11480 11336 11486 11348
rect 12069 11339 12127 11345
rect 12069 11336 12081 11339
rect 11480 11308 12081 11336
rect 11480 11296 11486 11308
rect 12069 11305 12081 11308
rect 12115 11305 12127 11339
rect 12069 11299 12127 11305
rect 11517 11271 11575 11277
rect 11517 11268 11529 11271
rect 11348 11240 11529 11268
rect 11517 11237 11529 11240
rect 11563 11237 11575 11271
rect 11517 11231 11575 11237
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 11664 11240 11928 11268
rect 11664 11228 11670 11240
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 11256 11200 11284 11228
rect 10735 11172 11284 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 11900 11209 11928 11240
rect 11974 11228 11980 11280
rect 12032 11268 12038 11280
rect 12345 11271 12403 11277
rect 12345 11268 12357 11271
rect 12032 11240 12357 11268
rect 12032 11228 12038 11240
rect 12345 11237 12357 11240
rect 12391 11237 12403 11271
rect 12345 11231 12403 11237
rect 11885 11203 11943 11209
rect 11532 11172 11744 11200
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 9272 11104 10609 11132
rect 9272 11092 9278 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 6114 11067 6172 11073
rect 6114 11033 6126 11067
rect 6160 11064 6172 11067
rect 6270 11064 6276 11076
rect 6160 11036 6276 11064
rect 6160 11033 6172 11036
rect 6114 11027 6172 11033
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 7282 11024 7288 11076
rect 7340 11024 7346 11076
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 8386 11064 8392 11076
rect 7432 11036 8392 11064
rect 7432 11024 7438 11036
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 10796 11064 10824 11095
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 11348 11064 11376 11160
rect 11422 11092 11428 11144
rect 11480 11132 11486 11144
rect 11532 11132 11560 11172
rect 11716 11141 11744 11172
rect 11885 11169 11897 11203
rect 11931 11169 11943 11203
rect 11885 11163 11943 11169
rect 11480 11104 11560 11132
rect 11609 11135 11667 11141
rect 11480 11092 11486 11104
rect 11609 11101 11621 11135
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 11839 11104 12020 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 10376 11036 11376 11064
rect 10376 11024 10382 11036
rect 11624 11008 11652 11095
rect 5902 10996 5908 11008
rect 4856 10968 5908 10996
rect 4856 10956 4862 10968
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6730 10996 6736 11008
rect 6052 10968 6736 10996
rect 6052 10956 6058 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 7745 10999 7803 11005
rect 7745 10965 7757 10999
rect 7791 10996 7803 10999
rect 7926 10996 7932 11008
rect 7791 10968 7932 10996
rect 7791 10965 7803 10968
rect 7745 10959 7803 10965
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 10962 10996 10968 11008
rect 8628 10968 10968 10996
rect 8628 10956 8634 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11606 10956 11612 11008
rect 11664 10956 11670 11008
rect 11992 10996 12020 11104
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 12667 11104 12756 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 12728 11008 12756 11104
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 12066 10996 12072 11008
rect 11992 10968 12072 10996
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 12526 10956 12532 11008
rect 12584 10956 12590 11008
rect 12710 10956 12716 11008
rect 12768 10956 12774 11008
rect 13170 10956 13176 11008
rect 13228 10956 13234 11008
rect 1104 10906 13984 10928
rect 1104 10854 4918 10906
rect 4970 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 5238 10906
rect 5290 10854 10918 10906
rect 10970 10854 10982 10906
rect 11034 10854 11046 10906
rect 11098 10854 11110 10906
rect 11162 10854 11174 10906
rect 11226 10854 11238 10906
rect 11290 10854 13984 10906
rect 1104 10832 13984 10854
rect 3602 10752 3608 10804
rect 3660 10752 3666 10804
rect 3887 10795 3945 10801
rect 3887 10761 3899 10795
rect 3933 10792 3945 10795
rect 3933 10764 4016 10792
rect 3933 10761 3945 10764
rect 3887 10755 3945 10761
rect 3988 10724 4016 10764
rect 4062 10752 4068 10804
rect 4120 10752 4126 10804
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4522 10792 4528 10804
rect 4479 10764 4528 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4893 10795 4951 10801
rect 4893 10761 4905 10795
rect 4939 10792 4951 10795
rect 4939 10764 5304 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 4338 10724 4344 10736
rect 3988 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10724 4402 10736
rect 4908 10724 4936 10755
rect 4396 10696 4936 10724
rect 4396 10684 4402 10696
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4154 10656 4160 10668
rect 4019 10628 4160 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4154 10616 4160 10628
rect 4212 10656 4218 10668
rect 4212 10628 4568 10656
rect 4212 10616 4218 10628
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4172 10560 4353 10588
rect 4172 10452 4200 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4540 10588 4568 10628
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4672 10628 4721 10656
rect 4672 10616 4678 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 4890 10656 4896 10668
rect 4847 10628 4896 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 4816 10588 4844 10619
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 4540 10560 4844 10588
rect 5169 10591 5227 10597
rect 4341 10551 4399 10557
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 5276 10588 5304 10764
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5408 10764 5457 10792
rect 5408 10752 5414 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 6420 10764 7297 10792
rect 6420 10752 6426 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 7374 10752 7380 10804
rect 7432 10752 7438 10804
rect 7466 10752 7472 10804
rect 7524 10752 7530 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 8076 10764 8585 10792
rect 8076 10752 8082 10764
rect 8573 10761 8585 10764
rect 8619 10792 8631 10795
rect 9766 10792 9772 10804
rect 8619 10764 9772 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 9766 10752 9772 10764
rect 9824 10792 9830 10804
rect 9824 10764 10180 10792
rect 9824 10752 9830 10764
rect 6457 10727 6515 10733
rect 6457 10724 6469 10727
rect 5736 10696 6469 10724
rect 5736 10668 5764 10696
rect 6457 10693 6469 10696
rect 6503 10693 6515 10727
rect 6457 10687 6515 10693
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 7392 10724 7420 10752
rect 6696 10696 7052 10724
rect 6696 10684 6702 10696
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 5994 10616 6000 10668
rect 6052 10616 6058 10668
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 6546 10656 6552 10668
rect 6227 10628 6552 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6546 10616 6552 10628
rect 6604 10656 6610 10668
rect 6822 10656 6828 10668
rect 6604 10628 6828 10656
rect 6604 10616 6610 10628
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7024 10665 7052 10696
rect 7300 10696 7420 10724
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7130 10659 7188 10665
rect 7130 10625 7142 10659
rect 7176 10656 7188 10659
rect 7300 10656 7328 10696
rect 7484 10665 7512 10752
rect 10042 10724 10048 10736
rect 9508 10696 10048 10724
rect 7176 10628 7328 10656
rect 7476 10659 7534 10665
rect 7176 10625 7188 10628
rect 7130 10619 7188 10625
rect 7476 10625 7488 10659
rect 7522 10625 7534 10659
rect 7476 10619 7534 10625
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7708 10628 7757 10656
rect 7708 10616 7714 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8352 10628 8401 10656
rect 8352 10616 8358 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 6012 10588 6040 10616
rect 5276 10560 6040 10588
rect 5169 10551 5227 10557
rect 4249 10523 4307 10529
rect 4249 10489 4261 10523
rect 4295 10520 4307 10523
rect 4798 10520 4804 10532
rect 4295 10492 4804 10520
rect 4295 10489 4307 10492
rect 4249 10483 4307 10489
rect 4798 10480 4804 10492
rect 4856 10520 4862 10532
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 4856 10492 5089 10520
rect 4856 10480 4862 10492
rect 5077 10489 5089 10492
rect 5123 10489 5135 10523
rect 5077 10483 5135 10489
rect 4614 10452 4620 10464
rect 4172 10424 4620 10452
rect 4614 10412 4620 10424
rect 4672 10452 4678 10464
rect 5184 10452 5212 10551
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7282 10588 7288 10600
rect 6963 10560 7288 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7340 10560 7573 10588
rect 7340 10548 7346 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 8404 10588 8432 10619
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8628 10628 8769 10656
rect 8628 10616 8634 10628
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9398 10656 9404 10668
rect 8996 10628 9404 10656
rect 8996 10616 9002 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 8956 10588 8984 10616
rect 8404 10560 8984 10588
rect 7561 10551 7619 10557
rect 5905 10523 5963 10529
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6362 10520 6368 10532
rect 5951 10492 6368 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6362 10480 6368 10492
rect 6420 10520 6426 10532
rect 6656 10520 6684 10548
rect 6420 10492 6684 10520
rect 9125 10523 9183 10529
rect 6420 10480 6426 10492
rect 9125 10489 9137 10523
rect 9171 10520 9183 10523
rect 9508 10520 9536 10696
rect 10042 10684 10048 10696
rect 10100 10684 10106 10736
rect 10152 10724 10180 10764
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11204 10764 11529 10792
rect 11204 10752 11210 10764
rect 11517 10761 11529 10764
rect 11563 10792 11575 10795
rect 12066 10792 12072 10804
rect 11563 10764 12072 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12216 10764 12633 10792
rect 12216 10752 12222 10764
rect 10152 10696 11192 10724
rect 10152 10665 10180 10696
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9692 10628 9873 10656
rect 9692 10532 9720 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10137 10659 10195 10665
rect 9999 10628 10088 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10060 10600 10088 10628
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10652 10628 10701 10656
rect 10652 10616 10658 10628
rect 10689 10625 10701 10628
rect 10735 10656 10747 10659
rect 10778 10656 10784 10668
rect 10735 10628 10784 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11054 10656 11060 10668
rect 11011 10628 11060 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11164 10656 11192 10696
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11675 10727 11733 10733
rect 11675 10724 11687 10727
rect 11296 10696 11687 10724
rect 11296 10684 11302 10696
rect 11675 10693 11687 10696
rect 11721 10693 11733 10727
rect 11675 10687 11733 10693
rect 11885 10727 11943 10733
rect 11885 10693 11897 10727
rect 11931 10693 11943 10727
rect 11885 10687 11943 10693
rect 11900 10656 11928 10687
rect 12268 10665 12296 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 13357 10727 13415 10733
rect 13357 10724 13369 10727
rect 12768 10696 13369 10724
rect 12768 10684 12774 10696
rect 13357 10693 13369 10696
rect 13403 10693 13415 10727
rect 13357 10687 13415 10693
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11164 10628 11989 10656
rect 11624 10600 11652 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10625 12311 10659
rect 12253 10619 12311 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 12986 10656 12992 10668
rect 12943 10628 12992 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 11606 10548 11612 10600
rect 11664 10548 11670 10600
rect 12176 10588 12204 10619
rect 12986 10616 12992 10628
rect 13044 10656 13050 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13044 10628 13553 10656
rect 13044 10616 13050 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13170 10588 13176 10600
rect 12176 10560 13176 10588
rect 9171 10492 9536 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 9582 10480 9588 10532
rect 9640 10480 9646 10532
rect 9674 10480 9680 10532
rect 9732 10480 9738 10532
rect 10778 10480 10784 10532
rect 10836 10480 10842 10532
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 11977 10523 12035 10529
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 12066 10520 12072 10532
rect 12023 10492 12072 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 4672 10424 5212 10452
rect 4672 10412 4678 10424
rect 5810 10412 5816 10464
rect 5868 10412 5874 10464
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6733 10455 6791 10461
rect 6733 10452 6745 10455
rect 6043 10424 6745 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6733 10421 6745 10424
rect 6779 10452 6791 10455
rect 6822 10452 6828 10464
rect 6779 10424 6828 10452
rect 6779 10421 6791 10424
rect 6733 10415 6791 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7742 10412 7748 10464
rect 7800 10412 7806 10464
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 10134 10452 10140 10464
rect 10091 10424 10140 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10376 10424 10517 10452
rect 10376 10412 10382 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10888 10452 10916 10483
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 12176 10464 12204 10560
rect 13170 10548 13176 10560
rect 13228 10588 13234 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 13228 10560 13277 10588
rect 13228 10548 13234 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 11146 10452 11152 10464
rect 10888 10424 11152 10452
rect 10505 10415 10563 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11480 10424 11713 10452
rect 11480 10412 11486 10424
rect 11701 10421 11713 10424
rect 11747 10452 11759 10455
rect 12158 10452 12164 10464
rect 11747 10424 12164 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 1104 10362 13984 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13984 10362
rect 1104 10288 13984 10310
rect 4249 10251 4307 10257
rect 4249 10217 4261 10251
rect 4295 10248 4307 10251
rect 4706 10248 4712 10260
rect 4295 10220 4712 10248
rect 4295 10217 4307 10220
rect 4249 10211 4307 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6641 10251 6699 10257
rect 6641 10248 6653 10251
rect 5868 10220 6653 10248
rect 5868 10208 5874 10220
rect 6641 10217 6653 10220
rect 6687 10217 6699 10251
rect 6641 10211 6699 10217
rect 4890 10140 4896 10192
rect 4948 10180 4954 10192
rect 6181 10183 6239 10189
rect 6181 10180 6193 10183
rect 4948 10152 6193 10180
rect 4948 10140 4954 10152
rect 6181 10149 6193 10152
rect 6227 10149 6239 10183
rect 6181 10143 6239 10149
rect 6457 10183 6515 10189
rect 6457 10149 6469 10183
rect 6503 10180 6515 10183
rect 6546 10180 6552 10192
rect 6503 10152 6552 10180
rect 6503 10149 6515 10152
rect 6457 10143 6515 10149
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 6656 10124 6684 10211
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7006 10248 7012 10260
rect 6880 10220 7012 10248
rect 6880 10208 6886 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7248 10220 7665 10248
rect 7248 10208 7254 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 7834 10208 7840 10260
rect 7892 10208 7898 10260
rect 8938 10208 8944 10260
rect 8996 10208 9002 10260
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9088 10220 10364 10248
rect 9088 10208 9094 10220
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 7469 10183 7527 10189
rect 7469 10180 7481 10183
rect 6788 10152 7481 10180
rect 6788 10140 6794 10152
rect 7469 10149 7481 10152
rect 7515 10149 7527 10183
rect 10336 10180 10364 10220
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 11756 10220 11897 10248
rect 11756 10208 11762 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 11885 10211 11943 10217
rect 12526 10180 12532 10192
rect 10336 10152 12532 10180
rect 7469 10143 7527 10149
rect 12526 10140 12532 10152
rect 12584 10180 12590 10192
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 12584 10152 12725 10180
rect 12584 10140 12590 10152
rect 12713 10149 12725 10152
rect 12759 10149 12771 10183
rect 12713 10143 12771 10149
rect 3881 10115 3939 10121
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 3927 10084 6500 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 6472 10056 6500 10084
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 6696 10084 7052 10112
rect 6696 10072 6702 10084
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6822 10044 6828 10056
rect 6595 10016 6828 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7024 10053 7052 10084
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7650 10112 7656 10124
rect 7248 10084 7656 10112
rect 7248 10072 7254 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 10321 10115 10379 10121
rect 7852 10084 8524 10112
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7374 10044 7380 10056
rect 7331 10016 7380 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7852 10044 7880 10084
rect 7524 10016 7880 10044
rect 7929 10047 7987 10053
rect 7524 10004 7530 10016
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8496 10044 8524 10084
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 11698 10112 11704 10124
rect 10367 10084 11704 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11790 10072 11796 10124
rect 11848 10072 11854 10124
rect 8570 10044 8576 10056
rect 8496 10016 8576 10044
rect 8021 10007 8079 10013
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 7834 9976 7840 9988
rect 6135 9948 7840 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4617 9911 4675 9917
rect 4617 9908 4629 9911
rect 4396 9880 4629 9908
rect 4396 9868 4402 9880
rect 4617 9877 4629 9880
rect 4663 9877 4675 9911
rect 4617 9871 4675 9877
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6420 9880 6837 9908
rect 6420 9868 6426 9880
rect 6825 9877 6837 9880
rect 6871 9877 6883 9911
rect 6825 9871 6883 9877
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 7944 9908 7972 10007
rect 8036 9976 8064 10007
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 10686 10044 10692 10056
rect 9646 10016 10692 10044
rect 8386 9976 8392 9988
rect 8036 9948 8392 9976
rect 8386 9936 8392 9948
rect 8444 9976 8450 9988
rect 9646 9976 9674 10016
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11808 10044 11836 10072
rect 11112 10016 11836 10044
rect 11112 10004 11118 10016
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12216 10016 12449 10044
rect 12216 10004 12222 10016
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 13044 10016 13093 10044
rect 13044 10004 13050 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 8444 9948 9674 9976
rect 8444 9936 8450 9948
rect 10042 9936 10048 9988
rect 10100 9985 10106 9988
rect 10100 9939 10112 9985
rect 10597 9979 10655 9985
rect 10597 9945 10609 9979
rect 10643 9945 10655 9979
rect 10695 9976 10723 10004
rect 12618 9976 12624 9988
rect 10695 9948 12624 9976
rect 10597 9939 10655 9945
rect 10100 9936 10106 9939
rect 7340 9880 7972 9908
rect 7340 9868 7346 9880
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 8536 9880 8677 9908
rect 8536 9868 8542 9880
rect 8665 9877 8677 9880
rect 8711 9908 8723 9911
rect 9030 9908 9036 9920
rect 8711 9880 9036 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 10612 9908 10640 9939
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 10686 9908 10692 9920
rect 9180 9880 10692 9908
rect 9180 9868 9186 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 12250 9908 12256 9920
rect 11296 9880 12256 9908
rect 11296 9868 11302 9880
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 1104 9818 13984 9840
rect 1104 9766 4918 9818
rect 4970 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 5238 9818
rect 5290 9766 10918 9818
rect 10970 9766 10982 9818
rect 11034 9766 11046 9818
rect 11098 9766 11110 9818
rect 11162 9766 11174 9818
rect 11226 9766 11238 9818
rect 11290 9766 13984 9818
rect 1104 9744 13984 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5077 9707 5135 9713
rect 5077 9704 5089 9707
rect 4856 9676 5089 9704
rect 4856 9664 4862 9676
rect 5077 9673 5089 9676
rect 5123 9673 5135 9707
rect 5077 9667 5135 9673
rect 6656 9676 7052 9704
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 4338 9636 4344 9648
rect 2832 9608 4344 9636
rect 2832 9596 2838 9608
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 5902 9636 5908 9648
rect 5276 9608 5908 9636
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3418 9568 3424 9580
rect 3283 9540 3424 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4154 9568 4160 9580
rect 3528 9540 4160 9568
rect 3528 9512 3556 9540
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 5276 9577 5304 9608
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 6656 9636 6684 9676
rect 6472 9608 6684 9636
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 6472 9568 6500 9608
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6788 9608 6837 9636
rect 6788 9596 6794 9608
rect 6825 9605 6837 9608
rect 6871 9636 6883 9639
rect 6917 9639 6975 9645
rect 6917 9636 6929 9639
rect 6871 9608 6929 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 6917 9605 6929 9608
rect 6963 9605 6975 9639
rect 7024 9636 7052 9676
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 9122 9704 9128 9716
rect 7892 9676 9128 9704
rect 7892 9664 7898 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9398 9664 9404 9716
rect 9456 9664 9462 9716
rect 10042 9664 10048 9716
rect 10100 9664 10106 9716
rect 10134 9664 10140 9716
rect 10192 9664 10198 9716
rect 10226 9664 10232 9716
rect 10284 9664 10290 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10560 9676 10916 9704
rect 10560 9664 10566 9676
rect 9416 9636 9444 9664
rect 7024 9608 7328 9636
rect 6917 9599 6975 9605
rect 5583 9540 6500 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 7300 9577 7328 9608
rect 9140 9608 9904 9636
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7331 9540 8984 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 2225 9503 2283 9509
rect 2225 9469 2237 9503
rect 2271 9500 2283 9503
rect 2958 9500 2964 9512
rect 2271 9472 2964 9500
rect 2271 9469 2283 9472
rect 2225 9463 2283 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3510 9500 3516 9512
rect 3375 9472 3516 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2639 9404 2881 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 3160 9432 3188 9463
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 5442 9460 5448 9512
rect 5500 9460 5506 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 6914 9500 6920 9512
rect 6779 9472 6920 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 3234 9432 3240 9444
rect 3160 9404 3240 9432
rect 2869 9395 2927 9401
rect 3234 9392 3240 9404
rect 3292 9432 3298 9444
rect 3896 9432 3924 9460
rect 7116 9444 7144 9531
rect 7098 9432 7104 9444
rect 3292 9404 3924 9432
rect 5552 9404 7104 9432
rect 3292 9392 3298 9404
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 3970 9364 3976 9376
rect 2731 9336 3976 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 5552 9373 5580 9404
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 8956 9376 8984 9540
rect 9030 9528 9036 9580
rect 9088 9528 9094 9580
rect 9140 9577 9168 9608
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 9140 9472 9321 9500
rect 9140 9444 9168 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9416 9500 9444 9531
rect 9582 9528 9588 9580
rect 9640 9528 9646 9580
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 9876 9500 9904 9608
rect 10152 9599 10180 9664
rect 10888 9636 10916 9676
rect 11698 9664 11704 9716
rect 11756 9664 11762 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 11885 9707 11943 9713
rect 11885 9704 11897 9707
rect 11848 9676 11897 9704
rect 11848 9664 11854 9676
rect 11885 9673 11897 9676
rect 11931 9673 11943 9707
rect 11885 9667 11943 9673
rect 10244 9608 10824 9636
rect 10888 9608 11008 9636
rect 10137 9593 10195 9599
rect 10137 9559 10149 9593
rect 10183 9559 10195 9593
rect 10137 9553 10195 9559
rect 10244 9500 10272 9608
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10796 9577 10824 9608
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10781 9571 10839 9577
rect 10643 9540 10732 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 9416 9472 9812 9500
rect 9876 9472 10272 9500
rect 9309 9463 9367 9469
rect 9784 9444 9812 9472
rect 9122 9392 9128 9444
rect 9180 9392 9186 9444
rect 9217 9435 9275 9441
rect 9217 9401 9229 9435
rect 9263 9432 9275 9435
rect 9674 9432 9680 9444
rect 9263 9404 9680 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9766 9392 9772 9444
rect 9824 9392 9830 9444
rect 10428 9432 10456 9528
rect 10704 9512 10732 9540
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10686 9460 10692 9512
rect 10744 9460 10750 9512
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 10980 9509 11008 9608
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 11296 9608 11529 9636
rect 11296 9596 11302 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11716 9636 11744 9664
rect 11716 9608 12112 9636
rect 11517 9599 11575 9605
rect 12084 9580 12112 9608
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9568 11207 9571
rect 11422 9568 11428 9580
rect 11195 9540 11428 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 11790 9568 11796 9580
rect 11747 9540 11796 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 12325 9571 12383 9577
rect 12325 9568 12337 9571
rect 12176 9540 12337 9568
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 12176 9500 12204 9540
rect 12325 9537 12337 9540
rect 12371 9537 12383 9571
rect 12325 9531 12383 9537
rect 11379 9472 12204 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 10152 9404 11008 9432
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6328 9336 6377 9364
rect 6328 9324 6334 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7374 9364 7380 9376
rect 6880 9336 7380 9364
rect 6880 9324 6886 9336
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 10152 9364 10180 9404
rect 10980 9376 11008 9404
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13412 9404 13461 9432
rect 13412 9392 13418 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 8996 9336 10180 9364
rect 8996 9324 9002 9336
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 10962 9324 10968 9376
rect 11020 9324 11026 9376
rect 1104 9274 13984 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13984 9274
rect 1104 9200 13984 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1578 9160 1584 9172
rect 1535 9132 1584 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2958 9120 2964 9172
rect 3016 9120 3022 9172
rect 3050 9120 3056 9172
rect 3108 9120 3114 9172
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 4246 9160 4252 9172
rect 3292 9132 4252 9160
rect 3292 9120 3298 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 6733 9163 6791 9169
rect 4672 9132 6684 9160
rect 4672 9120 4678 9132
rect 3068 9024 3096 9120
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 4706 9092 4712 9104
rect 3384 9064 4712 9092
rect 3384 9052 3390 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 3068 8996 3617 9024
rect 3605 8993 3617 8996
rect 3651 9024 3663 9027
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 3651 8996 4813 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2774 8956 2780 8968
rect 1728 8928 2780 8956
rect 1728 8916 1734 8928
rect 2774 8916 2780 8928
rect 2832 8956 2838 8968
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2832 8928 2881 8956
rect 2832 8916 2838 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 2602 8891 2660 8897
rect 2602 8888 2614 8891
rect 2004 8860 2614 8888
rect 2004 8848 2010 8860
rect 2602 8857 2614 8860
rect 2648 8857 2660 8891
rect 3160 8888 3188 8919
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 3878 8956 3884 8968
rect 3559 8928 3884 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 5000 8965 5028 9132
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 5810 9092 5816 9104
rect 5123 9064 5816 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 9024 5227 9027
rect 5442 9024 5448 9036
rect 5215 8996 5448 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 5442 8984 5448 8996
rect 5500 9024 5506 9036
rect 6656 9024 6684 9132
rect 6733 9129 6745 9163
rect 6779 9160 6791 9163
rect 7190 9160 7196 9172
rect 6779 9132 7196 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7466 9120 7472 9172
rect 7524 9120 7530 9172
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9769 9163 9827 9169
rect 9769 9160 9781 9163
rect 9640 9132 9781 9160
rect 9640 9120 9646 9132
rect 9769 9129 9781 9132
rect 9815 9129 9827 9163
rect 9769 9123 9827 9129
rect 9953 9163 10011 9169
rect 9953 9129 9965 9163
rect 9999 9129 10011 9163
rect 10410 9160 10416 9172
rect 9953 9123 10011 9129
rect 10060 9132 10416 9160
rect 7484 9024 7512 9120
rect 9416 9092 9444 9120
rect 9968 9092 9996 9123
rect 9416 9064 9996 9092
rect 9766 9024 9772 9036
rect 5500 8996 6500 9024
rect 5500 8984 5506 8996
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 3344 8888 3372 8916
rect 4522 8888 4528 8900
rect 3160 8860 3372 8888
rect 3712 8860 4528 8888
rect 2602 8851 2660 8857
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3234 8820 3240 8832
rect 2924 8792 3240 8820
rect 2924 8780 2930 8792
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3329 8823 3387 8829
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 3418 8820 3424 8832
rect 3375 8792 3424 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3418 8780 3424 8792
rect 3476 8820 3482 8832
rect 3712 8820 3740 8860
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 5276 8888 5304 8919
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5684 8928 5917 8956
rect 5684 8916 5690 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6472 8965 6500 8996
rect 6656 8996 7512 9024
rect 8864 8996 9772 9024
rect 6656 8965 6684 8996
rect 6840 8965 7052 8966
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6825 8959 7052 8965
rect 6825 8956 6837 8959
rect 6641 8919 6699 8925
rect 6748 8928 6837 8956
rect 6380 8888 6408 8916
rect 5276 8860 6408 8888
rect 3476 8792 3740 8820
rect 3476 8780 3482 8792
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 3936 8792 5549 8820
rect 3936 8780 3942 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 5537 8783 5595 8789
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6365 8823 6423 8829
rect 6365 8820 6377 8823
rect 6328 8792 6377 8820
rect 6328 8780 6334 8792
rect 6365 8789 6377 8792
rect 6411 8789 6423 8823
rect 6472 8820 6500 8919
rect 6546 8848 6552 8900
rect 6604 8888 6610 8900
rect 6748 8888 6776 8928
rect 6825 8925 6837 8928
rect 6871 8956 7052 8959
rect 8754 8956 8760 8968
rect 6871 8938 8760 8956
rect 6871 8925 6883 8938
rect 7024 8928 8760 8938
rect 6825 8919 6883 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 6604 8860 6776 8888
rect 6604 8848 6610 8860
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 8864 8888 8892 8996
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 10060 9033 10088 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 10928 9132 11253 9160
rect 10928 9120 10934 9132
rect 11241 9129 11253 9132
rect 11287 9129 11299 9163
rect 12710 9160 12716 9172
rect 11241 9123 11299 9129
rect 11532 9132 12716 9160
rect 11054 9052 11060 9104
rect 11112 9092 11118 9104
rect 11532 9092 11560 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 11112 9064 11560 9092
rect 11112 9052 11118 9064
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10652 8996 10824 9024
rect 10652 8984 10658 8996
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9858 8916 9864 8968
rect 9916 8950 9922 8968
rect 9953 8959 10011 8965
rect 9953 8950 9965 8959
rect 9916 8925 9965 8950
rect 9999 8925 10011 8959
rect 9916 8922 10011 8925
rect 9916 8916 9922 8922
rect 9953 8919 10011 8922
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 10796 8965 10824 8996
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10928 8996 11161 9024
rect 10928 8984 10934 8996
rect 11149 8993 11161 8996
rect 11195 9024 11207 9027
rect 11238 9024 11244 9036
rect 11195 8996 11244 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11388 8996 11468 9024
rect 11388 8984 11394 8996
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 6972 8860 8892 8888
rect 9140 8888 9168 8916
rect 9766 8888 9772 8900
rect 9140 8860 9772 8888
rect 6972 8848 6978 8860
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 10520 8888 10548 8919
rect 10428 8860 10548 8888
rect 6638 8820 6644 8832
rect 6472 8792 6644 8820
rect 6365 8783 6423 8789
rect 6638 8780 6644 8792
rect 6696 8820 6702 8832
rect 7742 8820 7748 8832
rect 6696 8792 7748 8820
rect 6696 8780 6702 8792
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10428 8820 10456 8860
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 9732 8792 10456 8820
rect 9732 8780 9738 8792
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10704 8820 10732 8919
rect 10962 8916 10968 8968
rect 11020 8916 11026 8968
rect 11440 8965 11468 8996
rect 11532 8965 11560 9064
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 11756 8996 11836 9024
rect 11756 8984 11762 8996
rect 11808 8965 11836 8996
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 11974 8956 11980 8968
rect 11931 8928 11980 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 11609 8891 11667 8897
rect 11609 8857 11621 8891
rect 11655 8857 11667 8891
rect 11609 8851 11667 8857
rect 10560 8792 10732 8820
rect 11624 8820 11652 8851
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 12314 8891 12372 8897
rect 12314 8888 12326 8891
rect 12216 8860 12326 8888
rect 12216 8848 12222 8860
rect 12314 8857 12326 8860
rect 12360 8857 12372 8891
rect 12314 8851 12372 8857
rect 12526 8848 12532 8900
rect 12584 8848 12590 8900
rect 12544 8820 12572 8848
rect 11624 8792 12572 8820
rect 10560 8780 10566 8792
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 13449 8823 13507 8829
rect 13449 8820 13461 8823
rect 13044 8792 13461 8820
rect 13044 8780 13050 8792
rect 13449 8789 13461 8792
rect 13495 8789 13507 8823
rect 13449 8783 13507 8789
rect 1104 8730 13984 8752
rect 1104 8678 4918 8730
rect 4970 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 5238 8730
rect 5290 8678 10918 8730
rect 10970 8678 10982 8730
rect 11034 8678 11046 8730
rect 11098 8678 11110 8730
rect 11162 8678 11174 8730
rect 11226 8678 11238 8730
rect 11290 8678 13984 8730
rect 1104 8656 13984 8678
rect 1946 8576 1952 8628
rect 2004 8576 2010 8628
rect 3970 8616 3976 8628
rect 2424 8588 3976 8616
rect 1596 8520 2360 8548
rect 1596 8492 1624 8520
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 2332 8489 2360 8520
rect 2424 8489 2452 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4157 8619 4215 8625
rect 4157 8616 4169 8619
rect 4080 8588 4169 8616
rect 3728 8551 3786 8557
rect 3728 8517 3740 8551
rect 3774 8548 3786 8551
rect 4080 8548 4108 8588
rect 4157 8585 4169 8588
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4304 8588 4445 8616
rect 4304 8576 4310 8588
rect 4433 8585 4445 8588
rect 4479 8616 4491 8619
rect 5810 8616 5816 8628
rect 4479 8588 5816 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6178 8576 6184 8628
rect 6236 8576 6242 8628
rect 6454 8616 6460 8628
rect 6288 8588 6460 8616
rect 6288 8560 6316 8588
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7558 8616 7564 8628
rect 7423 8588 7564 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 3774 8520 4108 8548
rect 3774 8517 3786 8520
rect 3728 8511 3786 8517
rect 4522 8508 4528 8560
rect 4580 8508 4586 8560
rect 6270 8508 6276 8560
rect 6328 8508 6334 8560
rect 6656 8548 6684 8576
rect 6472 8520 6684 8548
rect 6748 8548 6776 8579
rect 7558 8576 7564 8588
rect 7616 8616 7622 8628
rect 7616 8588 7788 8616
rect 7616 8576 7622 8588
rect 7760 8548 7788 8588
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 11422 8616 11428 8628
rect 8812 8588 11428 8616
rect 8812 8576 8818 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 12618 8576 12624 8628
rect 12676 8576 12682 8628
rect 9309 8551 9367 8557
rect 6748 8520 7512 8548
rect 7760 8520 8248 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 2832 8452 3985 8480
rect 2832 8440 2838 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 2130 8372 2136 8424
rect 2188 8372 2194 8424
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8381 2283 8415
rect 2866 8412 2872 8424
rect 2225 8375 2283 8381
rect 2516 8384 2872 8412
rect 2240 8344 2268 8375
rect 2516 8344 2544 8384
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 2240 8316 2544 8344
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 2958 8344 2964 8356
rect 2639 8316 2964 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 4172 8344 4200 8443
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 6472 8489 6500 8520
rect 5813 8483 5871 8489
rect 4672 8452 5396 8480
rect 4672 8440 4678 8452
rect 5368 8356 5396 8452
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 5859 8452 6469 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6914 8480 6920 8492
rect 6687 8452 6920 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7484 8489 7512 8520
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6564 8412 6592 8440
rect 5960 8384 6592 8412
rect 7208 8412 7236 8443
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 7760 8412 7788 8440
rect 7208 8384 7788 8412
rect 5960 8372 5966 8384
rect 5166 8344 5172 8356
rect 4172 8316 5172 8344
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5350 8304 5356 8356
rect 5408 8304 5414 8356
rect 5644 8344 5672 8372
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 5644 8316 7021 8344
rect 7009 8313 7021 8316
rect 7055 8313 7067 8347
rect 7009 8307 7067 8313
rect 4246 8236 4252 8288
rect 4304 8236 4310 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5718 8276 5724 8288
rect 5132 8248 5724 8276
rect 5132 8236 5138 8248
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8276 6055 8279
rect 6822 8276 6828 8288
rect 6043 8248 6828 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7098 8276 7104 8288
rect 6963 8248 7104 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 8220 8276 8248 8520
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 14090 8548 14096 8560
rect 9355 8520 14096 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9916 8452 10149 8480
rect 9916 8440 9922 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10502 8480 10508 8492
rect 10459 8452 10508 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 11146 8440 11152 8492
rect 11204 8440 11210 8492
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11606 8480 11612 8492
rect 11563 8452 11612 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12250 8480 12256 8492
rect 11931 8452 12256 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10796 8412 10824 8440
rect 9824 8384 10824 8412
rect 9824 8372 9830 8384
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10928 8384 11069 8412
rect 10928 8372 10934 8384
rect 11057 8381 11069 8384
rect 11103 8381 11115 8415
rect 11164 8412 11192 8440
rect 11716 8412 11744 8443
rect 11164 8384 11744 8412
rect 11057 8375 11115 8381
rect 10594 8304 10600 8356
rect 10652 8344 10658 8356
rect 11808 8344 11836 8443
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 12820 8412 12848 8443
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13372 8412 13400 8440
rect 12820 8384 13400 8412
rect 10652 8316 11836 8344
rect 10652 8304 10658 8316
rect 9766 8276 9772 8288
rect 8220 8248 9772 8276
rect 9766 8236 9772 8248
rect 9824 8276 9830 8288
rect 10226 8276 10232 8288
rect 9824 8248 10232 8276
rect 9824 8236 9830 8248
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 1104 8186 13984 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13984 8186
rect 1104 8112 13984 8134
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 4246 8072 4252 8084
rect 3375 8044 4252 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5074 8032 5080 8084
rect 5132 8032 5138 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 6365 8075 6423 8081
rect 6365 8072 6377 8075
rect 5408 8044 6377 8072
rect 5408 8032 5414 8044
rect 6365 8041 6377 8044
rect 6411 8041 6423 8075
rect 6365 8035 6423 8041
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 7190 8072 7196 8084
rect 6871 8044 7196 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7432 8044 8217 8072
rect 7432 8032 7438 8044
rect 8205 8041 8217 8044
rect 8251 8072 8263 8075
rect 8386 8072 8392 8084
rect 8251 8044 8392 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8496 8044 8953 8072
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3510 8004 3516 8016
rect 3099 7976 3516 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3510 7964 3516 7976
rect 3568 8004 3574 8016
rect 4062 8004 4068 8016
rect 3568 7976 4068 8004
rect 3568 7964 3574 7976
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4798 8004 4804 8016
rect 4212 7976 4804 8004
rect 4212 7964 4218 7976
rect 4798 7964 4804 7976
rect 4856 8004 4862 8016
rect 4985 8007 5043 8013
rect 4985 8004 4997 8007
rect 4856 7976 4997 8004
rect 4856 7964 4862 7976
rect 4985 7973 4997 7976
rect 5031 7973 5043 8007
rect 4985 7967 5043 7973
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 7742 8004 7748 8016
rect 5500 7976 7748 8004
rect 5500 7964 5506 7976
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 1670 7896 1676 7948
rect 1728 7896 1734 7948
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 4614 7936 4620 7948
rect 3476 7908 3556 7936
rect 3476 7896 3482 7908
rect 3528 7877 3556 7908
rect 3620 7908 4620 7936
rect 3620 7877 3648 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 6178 7896 6184 7948
rect 6236 7945 6242 7948
rect 6236 7939 6264 7945
rect 6252 7905 6264 7939
rect 6236 7899 6264 7905
rect 6236 7896 6242 7899
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6420 7908 6561 7936
rect 6420 7896 6426 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6696 7908 6929 7936
rect 6696 7896 6702 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 7374 7936 7380 7948
rect 7055 7908 7380 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 3513 7871 3571 7877
rect 3252 7840 3464 7868
rect 1940 7803 1998 7809
rect 1940 7769 1952 7803
rect 1986 7800 1998 7803
rect 3252 7800 3280 7840
rect 1986 7772 3280 7800
rect 3329 7803 3387 7809
rect 1986 7769 1998 7772
rect 1940 7763 1998 7769
rect 3329 7769 3341 7803
rect 3375 7769 3387 7803
rect 3436 7800 3464 7840
rect 3513 7837 3525 7871
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4706 7868 4712 7880
rect 4580 7840 4712 7868
rect 4580 7828 4586 7840
rect 4706 7828 4712 7840
rect 4764 7868 4770 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4764 7840 4813 7868
rect 4764 7828 4770 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 3786 7800 3792 7812
rect 3436 7772 3792 7800
rect 3329 7763 3387 7769
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 3344 7732 3372 7763
rect 3786 7760 3792 7772
rect 3844 7760 3850 7812
rect 4246 7760 4252 7812
rect 4304 7760 4310 7812
rect 5276 7800 5304 7831
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5442 7828 5448 7880
rect 5500 7862 5506 7880
rect 5537 7871 5595 7877
rect 5537 7862 5549 7871
rect 5500 7837 5549 7862
rect 5583 7837 5595 7871
rect 5500 7834 5595 7837
rect 5500 7828 5506 7834
rect 5537 7831 5595 7834
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5718 7828 5724 7880
rect 5776 7877 5782 7880
rect 5776 7868 5786 7877
rect 5776 7840 5821 7868
rect 5776 7831 5786 7840
rect 5776 7828 5782 7831
rect 5994 7828 6000 7880
rect 6052 7828 6058 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 8496 7877 8524 8044
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 8987 8044 9597 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9585 8041 9597 8044
rect 9631 8072 9643 8075
rect 10042 8072 10048 8084
rect 9631 8044 10048 8072
rect 9631 8041 9643 8044
rect 9585 8035 9643 8041
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 10594 8072 10600 8084
rect 10367 8044 10600 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10778 8072 10784 8084
rect 10735 8044 10784 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 9309 8007 9367 8013
rect 9309 8004 9321 8007
rect 8680 7976 9321 8004
rect 8680 7948 8708 7976
rect 9309 7973 9321 7976
rect 9355 8004 9367 8007
rect 9355 7976 9674 8004
rect 9355 7973 9367 7976
rect 9309 7967 9367 7973
rect 8662 7896 8668 7948
rect 8720 7896 8726 7948
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7156 7840 7297 7868
rect 7156 7828 7162 7840
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9171 7840 9505 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 5276 7772 8064 7800
rect 3602 7732 3608 7744
rect 3016 7704 3608 7732
rect 3016 7692 3022 7704
rect 3602 7692 3608 7704
rect 3660 7732 3666 7744
rect 4264 7732 4292 7760
rect 6012 7744 6040 7772
rect 3660 7704 4292 7732
rect 3660 7692 3666 7704
rect 5994 7692 6000 7744
rect 6052 7692 6058 7744
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 8036 7741 8064 7772
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 9140 7732 9168 7831
rect 9646 7800 9674 7976
rect 9766 7964 9772 8016
rect 9824 7964 9830 8016
rect 9784 7934 9812 7964
rect 9769 7928 9827 7934
rect 9769 7894 9781 7928
rect 9815 7894 9827 7928
rect 9769 7888 9827 7894
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10870 7868 10876 7880
rect 10827 7840 10876 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 10520 7800 10548 7828
rect 9646 7772 10548 7800
rect 8444 7704 9168 7732
rect 8444 7692 8450 7704
rect 9766 7692 9772 7744
rect 9824 7692 9830 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10796 7732 10824 7831
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 10100 7704 10824 7732
rect 10100 7692 10106 7704
rect 1104 7642 13984 7664
rect 1104 7590 4918 7642
rect 4970 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 5238 7642
rect 5290 7590 10918 7642
rect 10970 7590 10982 7642
rect 11034 7590 11046 7642
rect 11098 7590 11110 7642
rect 11162 7590 11174 7642
rect 11226 7590 11238 7642
rect 11290 7590 13984 7642
rect 1104 7568 13984 7590
rect 5534 7488 5540 7540
rect 5592 7488 5598 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6144 7500 6653 7528
rect 6144 7488 6150 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7558 7528 7564 7540
rect 6788 7500 7564 7528
rect 6788 7488 6794 7500
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 8662 7528 8668 7540
rect 8220 7500 8668 7528
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 7098 7460 7104 7472
rect 5408 7432 5948 7460
rect 5408 7420 5414 7432
rect 5920 7404 5948 7432
rect 6380 7432 7104 7460
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5684 7364 5733 7392
rect 5684 7352 5690 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5736 7268 5764 7355
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6380 7401 6408 7432
rect 7098 7420 7104 7432
rect 7156 7420 7162 7472
rect 6365 7395 6423 7401
rect 6052 7364 6094 7392
rect 6052 7352 6058 7364
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7392 7067 7395
rect 7282 7392 7288 7404
rect 7055 7364 7288 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 7524 7364 7573 7392
rect 7524 7352 7530 7364
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8220 7401 8248 7500
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 11572 7500 12434 7528
rect 11572 7488 11578 7500
rect 8386 7420 8392 7472
rect 8444 7420 8450 7472
rect 8507 7463 8565 7469
rect 8507 7429 8519 7463
rect 8553 7460 8565 7463
rect 8553 7432 8800 7460
rect 8553 7429 8565 7432
rect 8507 7423 8565 7429
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7800 7364 8033 7392
rect 7800 7352 7806 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 6454 7284 6460 7336
rect 6512 7284 6518 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6730 7324 6736 7336
rect 6687 7296 6736 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7392 7324 7420 7352
rect 7650 7324 7656 7336
rect 7392 7296 7656 7324
rect 7650 7284 7656 7296
rect 7708 7324 7714 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7708 7296 8677 7324
rect 7708 7284 7714 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 5718 7216 5724 7268
rect 5776 7256 5782 7268
rect 5776 7228 6960 7256
rect 5776 7216 5782 7228
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6454 7188 6460 7200
rect 5868 7160 6460 7188
rect 5868 7148 5874 7160
rect 6454 7148 6460 7160
rect 6512 7188 6518 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6512 7160 6837 7188
rect 6512 7148 6518 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6932 7188 6960 7228
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 8772 7256 8800 7432
rect 10704 7432 11744 7460
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 10704 7401 10732 7432
rect 11716 7404 11744 7432
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 9968 7364 10701 7392
rect 9968 7256 9996 7364
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11422 7392 11428 7404
rect 10919 7364 11428 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12406 7401 12434 7500
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11940 7364 11989 7392
rect 11940 7352 11946 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12353 7395 12434 7401
rect 12353 7361 12365 7395
rect 12399 7364 12434 7395
rect 12399 7361 12411 7364
rect 12353 7355 12411 7361
rect 11514 7324 11520 7336
rect 8628 7228 9996 7256
rect 10060 7296 11520 7324
rect 8628 7216 8634 7228
rect 10060 7200 10088 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 11992 7324 12020 7355
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 11992 7296 12449 7324
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 10042 7188 10048 7200
rect 6932 7160 10048 7188
rect 6825 7151 6883 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10284 7160 10701 7188
rect 10284 7148 10290 7160
rect 10689 7157 10701 7160
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 1104 7098 13984 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13984 7098
rect 1104 7024 13984 7046
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6273 6987 6331 6993
rect 6273 6984 6285 6987
rect 5960 6956 6285 6984
rect 5960 6944 5966 6956
rect 6273 6953 6285 6956
rect 6319 6953 6331 6987
rect 6273 6947 6331 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7742 6984 7748 6996
rect 7248 6956 7748 6984
rect 7248 6944 7254 6956
rect 7742 6944 7748 6956
rect 7800 6984 7806 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7800 6956 7941 6984
rect 7800 6944 7806 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 9030 6984 9036 6996
rect 7929 6947 7987 6953
rect 8588 6956 9036 6984
rect 6089 6919 6147 6925
rect 6089 6885 6101 6919
rect 6135 6885 6147 6919
rect 6089 6879 6147 6885
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 3970 6848 3976 6860
rect 2924 6820 3976 6848
rect 2924 6808 2930 6820
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 6104 6848 6132 6879
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 7340 6888 7573 6916
rect 7340 6876 7346 6888
rect 7561 6885 7573 6888
rect 7607 6885 7619 6919
rect 7561 6879 7619 6885
rect 7466 6848 7472 6860
rect 6104 6820 7472 6848
rect 7466 6808 7472 6820
rect 7524 6848 7530 6860
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7524 6820 7849 6848
rect 7524 6808 7530 6820
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 7944 6848 7972 6947
rect 8588 6848 8616 6956
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 9585 6987 9643 6993
rect 9585 6984 9597 6987
rect 9548 6956 9597 6984
rect 9548 6944 9554 6956
rect 9585 6953 9597 6956
rect 9631 6953 9643 6987
rect 9585 6947 9643 6953
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10505 6987 10563 6993
rect 10505 6984 10517 6987
rect 9916 6956 10517 6984
rect 9916 6944 9922 6956
rect 10505 6953 10517 6956
rect 10551 6953 10563 6987
rect 10505 6947 10563 6953
rect 8662 6876 8668 6928
rect 8720 6876 8726 6928
rect 9950 6876 9956 6928
rect 10008 6876 10014 6928
rect 11333 6919 11391 6925
rect 11333 6885 11345 6919
rect 11379 6885 11391 6919
rect 11333 6879 11391 6885
rect 7944 6820 8616 6848
rect 7837 6811 7895 6817
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 2958 6672 2964 6724
rect 3016 6712 3022 6724
rect 4724 6712 4752 6743
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 4965 6783 5023 6789
rect 4965 6780 4977 6783
rect 4856 6752 4977 6780
rect 4856 6740 4862 6752
rect 4965 6749 4977 6752
rect 5011 6749 5023 6783
rect 4965 6743 5023 6749
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6914 6780 6920 6792
rect 6503 6752 6920 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6914 6740 6920 6752
rect 6972 6780 6978 6792
rect 7098 6780 7104 6792
rect 6972 6752 7104 6780
rect 6972 6740 6978 6752
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 3016 6684 4844 6712
rect 3016 6672 3022 6684
rect 4816 6656 4844 6684
rect 3234 6604 3240 6656
rect 3292 6604 3298 6656
rect 4798 6604 4804 6656
rect 4856 6604 4862 6656
rect 7852 6644 7880 6811
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8588 6789 8616 6820
rect 8680 6848 8708 6876
rect 10045 6851 10103 6857
rect 8680 6820 9720 6848
rect 8680 6789 8708 6820
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 8404 6712 8432 6743
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 8812 6752 9260 6780
rect 8812 6740 8818 6752
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 8076 6684 8953 6712
rect 8076 6672 8082 6684
rect 8941 6681 8953 6684
rect 8987 6712 8999 6715
rect 9122 6712 9128 6724
rect 8987 6684 9128 6712
rect 8987 6681 8999 6684
rect 8941 6675 8999 6681
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 9232 6712 9260 6752
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9692 6780 9720 6820
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 10226 6848 10232 6860
rect 10091 6820 10232 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 11348 6848 11376 6879
rect 10428 6820 11376 6848
rect 11517 6851 11575 6857
rect 10428 6789 10456 6820
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11563 6820 11989 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 9692 6752 10425 6780
rect 9401 6743 9459 6749
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 9416 6712 9444 6743
rect 9232 6684 9444 6712
rect 9674 6672 9680 6724
rect 9732 6672 9738 6724
rect 9766 6672 9772 6724
rect 9824 6672 9830 6724
rect 10134 6672 10140 6724
rect 10192 6672 10198 6724
rect 8754 6644 8760 6656
rect 7852 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 10704 6644 10732 6743
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 11606 6780 11612 6792
rect 10836 6752 11612 6780
rect 10836 6740 10842 6752
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 11793 6783 11851 6789
rect 11793 6780 11805 6783
rect 11756 6752 11805 6780
rect 11756 6740 11762 6752
rect 11793 6749 11805 6752
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6780 12219 6783
rect 13446 6780 13452 6792
rect 12207 6752 13452 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6712 11115 6715
rect 11330 6712 11336 6724
rect 11103 6684 11336 6712
rect 11103 6681 11115 6684
rect 11057 6675 11115 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 9364 6616 10732 6644
rect 9364 6604 9370 6616
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 10965 6647 11023 6653
rect 10965 6644 10977 6647
rect 10836 6616 10977 6644
rect 10836 6604 10842 6616
rect 10965 6613 10977 6616
rect 11011 6613 11023 6647
rect 10965 6607 11023 6613
rect 12342 6604 12348 6656
rect 12400 6604 12406 6656
rect 1104 6554 13984 6576
rect 1104 6502 4918 6554
rect 4970 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 5238 6554
rect 5290 6502 10918 6554
rect 10970 6502 10982 6554
rect 11034 6502 11046 6554
rect 11098 6502 11110 6554
rect 11162 6502 11174 6554
rect 11226 6502 11238 6554
rect 11290 6502 13984 6554
rect 1104 6480 13984 6502
rect 3050 6400 3056 6452
rect 3108 6400 3114 6452
rect 3234 6400 3240 6452
rect 3292 6400 3298 6452
rect 3786 6440 3792 6452
rect 3620 6412 3792 6440
rect 2613 6307 2671 6313
rect 2613 6273 2625 6307
rect 2659 6304 2671 6307
rect 2869 6307 2927 6313
rect 2659 6276 2820 6304
rect 2659 6273 2671 6276
rect 2613 6267 2671 6273
rect 2792 6236 2820 6276
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 2958 6304 2964 6316
rect 2915 6276 2964 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 2792 6208 3004 6236
rect 2976 6177 3004 6208
rect 2961 6171 3019 6177
rect 2961 6137 2973 6171
rect 3007 6137 3019 6171
rect 3068 6168 3096 6400
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3252 6304 3280 6400
rect 3620 6381 3648 6412
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 8938 6440 8944 6452
rect 6328 6412 8944 6440
rect 6328 6400 6334 6412
rect 8938 6400 8944 6412
rect 8996 6440 9002 6452
rect 10042 6440 10048 6452
rect 8996 6412 10048 6440
rect 8996 6400 9002 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11330 6440 11336 6452
rect 10980 6412 11336 6440
rect 3513 6375 3571 6381
rect 3513 6341 3525 6375
rect 3559 6341 3571 6375
rect 3513 6335 3571 6341
rect 3605 6375 3663 6381
rect 3605 6341 3617 6375
rect 3651 6341 3663 6375
rect 6914 6372 6920 6384
rect 3605 6335 3663 6341
rect 3712 6344 6920 6372
rect 3191 6276 3280 6304
rect 3421 6307 3479 6313
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3528 6304 3556 6335
rect 3712 6304 3740 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7300 6344 7512 6372
rect 3528 6276 3740 6304
rect 3789 6307 3847 6313
rect 3421 6267 3479 6273
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 3436 6236 3464 6267
rect 3436 6208 3648 6236
rect 3620 6180 3648 6208
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 3068 6140 3249 6168
rect 2961 6131 3019 6137
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 3602 6128 3608 6180
rect 3660 6128 3666 6180
rect 1489 6103 1547 6109
rect 1489 6069 1501 6103
rect 1535 6100 1547 6103
rect 1670 6100 1676 6112
rect 1535 6072 1676 6100
rect 1535 6069 1547 6072
rect 1489 6063 1547 6069
rect 1670 6060 1676 6072
rect 1728 6100 1734 6112
rect 3804 6100 3832 6267
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4062 6264 4068 6316
rect 4120 6264 4126 6316
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6304 7251 6307
rect 7300 6304 7328 6344
rect 7484 6316 7512 6344
rect 7760 6344 8340 6372
rect 7239 6276 7328 6304
rect 7239 6273 7251 6276
rect 7193 6267 7251 6273
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 7760 6313 7788 6344
rect 8312 6316 8340 6344
rect 8570 6332 8576 6384
rect 8628 6332 8634 6384
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9214 6372 9220 6384
rect 9088 6344 9220 6372
rect 9088 6332 9094 6344
rect 9214 6332 9220 6344
rect 9272 6372 9278 6384
rect 9272 6344 9845 6372
rect 9272 6332 9278 6344
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7524 6276 7573 6304
rect 7524 6264 7530 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9582 6304 9588 6316
rect 8812 6276 9588 6304
rect 8812 6264 8818 6276
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9817 6304 9845 6344
rect 10980 6316 11008 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 11480 6344 11529 6372
rect 11480 6332 11486 6344
rect 11517 6341 11529 6344
rect 11563 6341 11575 6375
rect 11517 6335 11575 6341
rect 9817 6276 9904 6304
rect 3988 6236 4016 6264
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 3988 6208 4261 6236
rect 4249 6205 4261 6208
rect 4295 6236 4307 6239
rect 4706 6236 4712 6248
rect 4295 6208 4712 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 8478 6236 8484 6248
rect 6757 6208 8484 6236
rect 4522 6128 4528 6180
rect 4580 6168 4586 6180
rect 6757 6168 6785 6208
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8772 6236 8800 6264
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8772 6208 8953 6236
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9030 6196 9036 6248
rect 9088 6196 9094 6248
rect 9876 6236 9904 6276
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10781 6307 10839 6313
rect 10183 6276 10272 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10244 6236 10272 6276
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10962 6304 10968 6316
rect 10827 6276 10968 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11330 6304 11336 6316
rect 11287 6276 11336 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 9232 6208 9845 6236
rect 9876 6208 10272 6236
rect 13265 6239 13323 6245
rect 4580 6140 6785 6168
rect 4580 6128 4586 6140
rect 7650 6128 7656 6180
rect 7708 6128 7714 6180
rect 1728 6072 3832 6100
rect 1728 6060 1734 6072
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 4614 6100 4620 6112
rect 4479 6072 4620 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 7098 6060 7104 6112
rect 7156 6060 7162 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8478 6100 8484 6112
rect 8352 6072 8484 6100
rect 8352 6060 8358 6072
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9048 6109 9076 6196
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9232 6168 9260 6208
rect 9180 6140 9260 6168
rect 9180 6128 9186 6140
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 9493 6171 9551 6177
rect 9493 6168 9505 6171
rect 9364 6140 9505 6168
rect 9364 6128 9370 6140
rect 9493 6137 9505 6140
rect 9539 6137 9551 6171
rect 9817 6168 9845 6208
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13354 6236 13360 6248
rect 13311 6208 13360 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 9493 6131 9551 6137
rect 9600 6140 9720 6168
rect 9817 6140 9996 6168
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 9600 6100 9628 6140
rect 9456 6072 9628 6100
rect 9692 6100 9720 6140
rect 9766 6100 9772 6112
rect 9692 6072 9772 6100
rect 9456 6060 9462 6072
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9968 6100 9996 6140
rect 10962 6100 10968 6112
rect 9968 6072 10968 6100
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 1104 6010 13984 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13984 6010
rect 1104 5936 13984 5958
rect 2958 5896 2964 5908
rect 2240 5868 2964 5896
rect 2240 5769 2268 5868
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3878 5896 3884 5908
rect 3384 5868 3884 5896
rect 3384 5856 3390 5868
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4341 5899 4399 5905
rect 4341 5896 4353 5899
rect 4120 5868 4353 5896
rect 4120 5856 4126 5868
rect 4341 5865 4353 5868
rect 4387 5865 4399 5899
rect 4341 5859 4399 5865
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 7432 5868 8125 5896
rect 7432 5856 7438 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8444 5868 8677 5896
rect 8444 5856 8450 5868
rect 8665 5865 8677 5868
rect 8711 5896 8723 5899
rect 9769 5899 9827 5905
rect 9769 5896 9781 5899
rect 8711 5868 9781 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 9769 5865 9781 5868
rect 9815 5865 9827 5899
rect 9769 5859 9827 5865
rect 10134 5856 10140 5908
rect 10192 5856 10198 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11020 5868 11713 5896
rect 11020 5856 11026 5868
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 11701 5859 11759 5865
rect 4430 5828 4436 5840
rect 3436 5800 4436 5828
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2240 5692 2268 5723
rect 2314 5692 2320 5704
rect 2240 5664 2320 5692
rect 2133 5655 2191 5661
rect 2148 5624 2176 5655
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 3436 5692 3464 5800
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7800 5800 7849 5828
rect 7800 5788 7806 5800
rect 7837 5797 7849 5800
rect 7883 5797 7895 5831
rect 9122 5828 9128 5840
rect 7837 5791 7895 5797
rect 8312 5800 9128 5828
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 3970 5760 3976 5772
rect 3660 5732 3976 5760
rect 3660 5720 3666 5732
rect 3970 5720 3976 5732
rect 4028 5760 4034 5772
rect 6457 5763 6515 5769
rect 6457 5760 6469 5763
rect 4028 5732 4200 5760
rect 4028 5720 4034 5732
rect 4172 5701 4200 5732
rect 5644 5732 6469 5760
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2424 5664 3464 5692
rect 3620 5664 3801 5692
rect 2424 5624 2452 5664
rect 2148 5596 2452 5624
rect 2492 5627 2550 5633
rect 2492 5593 2504 5627
rect 2538 5624 2550 5627
rect 2958 5624 2964 5636
rect 2538 5596 2964 5624
rect 2538 5593 2550 5596
rect 2492 5587 2550 5593
rect 2958 5584 2964 5596
rect 3016 5584 3022 5636
rect 3620 5568 3648 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3789 5655 3847 5661
rect 3896 5664 4077 5692
rect 3694 5584 3700 5636
rect 3752 5624 3758 5636
rect 3896 5624 3924 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 3752 5596 3924 5624
rect 3973 5627 4031 5633
rect 3752 5584 3758 5596
rect 3973 5593 3985 5627
rect 4019 5593 4031 5627
rect 3973 5587 4031 5593
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1820 5528 1961 5556
rect 1820 5516 1826 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 1949 5519 2007 5525
rect 3602 5516 3608 5568
rect 3660 5516 3666 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 3988 5556 4016 5587
rect 5644 5568 5672 5732
rect 6457 5729 6469 5732
rect 6503 5729 6515 5763
rect 7852 5760 7880 5791
rect 8312 5772 8340 5800
rect 9122 5788 9128 5800
rect 9180 5788 9186 5840
rect 9582 5788 9588 5840
rect 9640 5828 9646 5840
rect 9640 5800 9904 5828
rect 9640 5788 9646 5800
rect 7852 5732 8248 5760
rect 6457 5723 6515 5729
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 7834 5692 7840 5704
rect 6411 5664 7840 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8220 5701 8248 5732
rect 8294 5720 8300 5772
rect 8352 5720 8358 5772
rect 9674 5760 9680 5772
rect 8956 5732 9680 5760
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8956 5703 8984 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9876 5769 9904 5800
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 8941 5697 8999 5703
rect 8536 5664 8892 5692
rect 8536 5652 8542 5664
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 6702 5627 6760 5633
rect 6702 5624 6714 5627
rect 6604 5596 6714 5624
rect 6604 5584 6610 5596
rect 6702 5593 6714 5596
rect 6748 5593 6760 5627
rect 8864 5624 8892 5664
rect 8941 5663 8953 5697
rect 8987 5663 8999 5697
rect 8941 5657 8999 5663
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 9088 5664 9137 5692
rect 9088 5652 9094 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9214 5652 9220 5704
rect 9272 5652 9278 5704
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9600 5664 9781 5692
rect 9324 5624 9352 5652
rect 8864 5596 9352 5624
rect 6702 5587 6760 5593
rect 3936 5528 4016 5556
rect 3936 5516 3942 5528
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 4856 5528 5089 5556
rect 4856 5516 4862 5528
rect 5077 5525 5089 5528
rect 5123 5556 5135 5559
rect 5626 5556 5632 5568
rect 5123 5528 5632 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9600 5556 9628 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 9364 5528 9628 5556
rect 9364 5516 9370 5528
rect 9674 5516 9680 5568
rect 9732 5516 9738 5568
rect 10060 5556 10088 5652
rect 10152 5624 10180 5856
rect 12066 5788 12072 5840
rect 12124 5788 12130 5840
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 12158 5692 12164 5704
rect 10367 5664 12164 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 12158 5652 12164 5664
rect 12216 5692 12222 5704
rect 13354 5692 13360 5704
rect 12216 5664 13360 5692
rect 12216 5652 12222 5664
rect 13354 5652 13360 5664
rect 13412 5692 13418 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 13412 5664 13461 5692
rect 13412 5652 13418 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 10566 5627 10624 5633
rect 10566 5624 10578 5627
rect 10152 5596 10578 5624
rect 10566 5593 10578 5596
rect 10612 5593 10624 5627
rect 10566 5587 10624 5593
rect 13170 5584 13176 5636
rect 13228 5633 13234 5636
rect 13228 5587 13240 5633
rect 13228 5584 13234 5587
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 10060 5528 10149 5556
rect 10137 5525 10149 5528
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 1104 5466 13984 5488
rect 1104 5414 4918 5466
rect 4970 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 5238 5466
rect 5290 5414 10918 5466
rect 10970 5414 10982 5466
rect 11034 5414 11046 5466
rect 11098 5414 11110 5466
rect 11162 5414 11174 5466
rect 11226 5414 11238 5466
rect 11290 5414 13984 5466
rect 1104 5392 13984 5414
rect 2958 5312 2964 5364
rect 3016 5312 3022 5364
rect 3326 5312 3332 5364
rect 3384 5312 3390 5364
rect 3878 5352 3884 5364
rect 3436 5324 3884 5352
rect 3344 5284 3372 5312
rect 3436 5293 3464 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 4430 5312 4436 5364
rect 4488 5312 4494 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4724 5324 5089 5352
rect 1504 5256 2360 5284
rect 1504 5225 1532 5256
rect 2332 5228 2360 5256
rect 3160 5256 3372 5284
rect 3421 5287 3479 5293
rect 1762 5225 1768 5228
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5185 1547 5219
rect 1756 5216 1768 5225
rect 1723 5188 1768 5216
rect 1489 5179 1547 5185
rect 1756 5179 1768 5188
rect 1762 5176 1768 5179
rect 1820 5176 1826 5228
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 3160 5225 3188 5256
rect 3421 5253 3433 5287
rect 3467 5253 3479 5287
rect 3421 5247 3479 5253
rect 3513 5287 3571 5293
rect 3513 5253 3525 5287
rect 3559 5284 3571 5287
rect 4522 5284 4528 5296
rect 3559 5256 4528 5284
rect 3559 5253 3571 5256
rect 3513 5247 3571 5253
rect 4522 5244 4528 5256
rect 4580 5244 4586 5296
rect 4724 5228 4752 5324
rect 5077 5321 5089 5324
rect 5123 5352 5135 5355
rect 7374 5352 7380 5364
rect 5123 5324 7380 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5352 7711 5355
rect 9030 5352 9036 5364
rect 7699 5324 9036 5352
rect 7699 5321 7711 5324
rect 7653 5315 7711 5321
rect 6365 5287 6423 5293
rect 6365 5253 6377 5287
rect 6411 5284 6423 5287
rect 6914 5284 6920 5296
rect 6411 5256 6920 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 7668 5284 7696 5315
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 9456 5324 10425 5352
rect 9456 5312 9462 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 10889 5355 10947 5361
rect 10889 5352 10901 5355
rect 10836 5324 10901 5352
rect 10836 5312 10842 5324
rect 10889 5321 10901 5324
rect 10935 5321 10947 5355
rect 10889 5315 10947 5321
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11848 5324 11897 5352
rect 11848 5312 11854 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 13446 5312 13452 5364
rect 13504 5312 13510 5364
rect 7024 5256 7696 5284
rect 7837 5287 7895 5293
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3970 5216 3976 5228
rect 3651 5188 3976 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3252 5148 3280 5179
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 2884 5120 3280 5148
rect 2884 5024 2912 5120
rect 3789 5083 3847 5089
rect 3789 5049 3801 5083
rect 3835 5080 3847 5083
rect 4632 5080 4660 5179
rect 4706 5176 4712 5228
rect 4764 5176 4770 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 3835 5052 4660 5080
rect 3835 5049 3847 5052
rect 3789 5043 3847 5049
rect 4706 5040 4712 5092
rect 4764 5080 4770 5092
rect 4908 5080 4936 5179
rect 5534 5176 5540 5228
rect 5592 5220 5598 5228
rect 5592 5192 5662 5220
rect 5592 5176 5598 5192
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5634 5148 5662 5192
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6512 5188 6561 5216
rect 6512 5176 6518 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 7024 5225 7052 5256
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8294 5284 8300 5296
rect 7883 5256 8300 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8386 5244 8392 5296
rect 8444 5284 8450 5296
rect 8941 5287 8999 5293
rect 8941 5284 8953 5287
rect 8444 5256 8953 5284
rect 8444 5244 8450 5256
rect 8941 5253 8953 5256
rect 8987 5253 8999 5287
rect 8941 5247 8999 5253
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7156 5188 7297 5216
rect 7156 5176 7162 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8312 5216 8340 5244
rect 8159 5188 8340 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 5634 5120 6837 5148
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 5718 5080 5724 5092
rect 4764 5052 5724 5080
rect 4764 5040 4770 5052
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 6365 5083 6423 5089
rect 6365 5049 6377 5083
rect 6411 5080 6423 5083
rect 6546 5080 6552 5092
rect 6411 5052 6552 5080
rect 6411 5049 6423 5052
rect 6365 5043 6423 5049
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 7300 5080 7328 5179
rect 8036 5148 8064 5179
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8496 5148 8524 5176
rect 8036 5120 8524 5148
rect 8772 5080 8800 5179
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9416 5225 9444 5312
rect 9490 5244 9496 5296
rect 9548 5284 9554 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 9548 5256 10701 5284
rect 9548 5244 9554 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 11532 5284 11560 5312
rect 12342 5293 12348 5296
rect 12336 5284 12348 5293
rect 11532 5256 12020 5284
rect 12303 5256 12348 5284
rect 10689 5247 10747 5253
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 9180 5188 9229 5216
rect 9180 5176 9186 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9858 5176 9864 5228
rect 9916 5176 9922 5228
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10226 5216 10232 5228
rect 10091 5188 10232 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11330 5216 11336 5228
rect 10643 5188 11336 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11992 5225 12020 5256
rect 12336 5247 12348 5256
rect 12342 5244 12348 5247
rect 12400 5244 12406 5296
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5216 12127 5219
rect 12158 5216 12164 5228
rect 12115 5188 12164 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 7300 5052 8800 5080
rect 10888 5052 11529 5080
rect 2866 4972 2872 5024
rect 2924 4972 2930 5024
rect 8312 5021 8340 5052
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 4981 8355 5015
rect 8297 4975 8355 4981
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 9122 4972 9128 5024
rect 9180 4972 9186 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9364 4984 9413 5012
rect 9364 4972 9370 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 10042 4972 10048 5024
rect 10100 4972 10106 5024
rect 10888 5021 10916 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 10873 5015 10931 5021
rect 10873 4981 10885 5015
rect 10919 4981 10931 5015
rect 10873 4975 10931 4981
rect 11054 4972 11060 5024
rect 11112 4972 11118 5024
rect 1104 4922 13984 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13984 4922
rect 1104 4848 13984 4870
rect 6638 4768 6644 4820
rect 6696 4768 6702 4820
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 9490 4808 9496 4820
rect 6788 4780 9496 4808
rect 6788 4768 6794 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10686 4808 10692 4820
rect 9600 4780 10692 4808
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4641 4215 4675
rect 4157 4635 4215 4641
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3476 4576 3985 4604
rect 3476 4564 3482 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 4172 4604 4200 4635
rect 4706 4604 4712 4616
rect 4172 4576 4712 4604
rect 3973 4567 4031 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4856 4576 4997 4604
rect 4856 4564 4862 4576
rect 4985 4573 4997 4576
rect 5031 4573 5043 4607
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4985 4567 5043 4573
rect 5092 4576 5273 4604
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 5092 4536 5120 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 5534 4604 5540 4616
rect 5399 4576 5540 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 6656 4604 6684 4768
rect 9600 4740 9628 4780
rect 7392 4712 9628 4740
rect 7392 4684 7420 4712
rect 9674 4700 9680 4752
rect 9732 4700 9738 4752
rect 9769 4743 9827 4749
rect 9769 4709 9781 4743
rect 9815 4740 9827 4743
rect 9950 4740 9956 4752
rect 9815 4712 9956 4740
rect 9815 4709 9827 4712
rect 9769 4703 9827 4709
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 8386 4672 8392 4684
rect 8220 4644 8392 4672
rect 8220 4613 8248 4644
rect 8386 4632 8392 4644
rect 8444 4672 8450 4684
rect 9122 4672 9128 4684
rect 8444 4644 9128 4672
rect 8444 4632 8450 4644
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9692 4672 9720 4700
rect 10152 4681 10180 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11054 4768 11060 4820
rect 11112 4768 11118 4820
rect 10137 4675 10195 4681
rect 9508 4644 9996 4672
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 6656 4576 8217 4604
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8570 4604 8576 4616
rect 8343 4576 8576 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8570 4564 8576 4576
rect 8628 4604 8634 4616
rect 9306 4604 9312 4616
rect 8628 4576 9312 4604
rect 8628 4564 8634 4576
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9508 4613 9536 4644
rect 9968 4613 9996 4644
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4573 9551 4607
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9493 4567 9551 4573
rect 9646 4576 9873 4604
rect 4212 4508 5120 4536
rect 5169 4539 5227 4545
rect 4212 4496 4218 4508
rect 5169 4505 5181 4539
rect 5215 4505 5227 4539
rect 5736 4536 5764 4564
rect 9646 4548 9674 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4573 10011 4607
rect 11072 4604 11100 4768
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 11072 4576 11161 4604
rect 9953 4567 10011 4573
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 6730 4536 6736 4548
rect 5736 4508 6736 4536
rect 5169 4499 5227 4505
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 5184 4468 5212 4499
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 8128 4508 8432 4536
rect 8128 4480 8156 4508
rect 5350 4468 5356 4480
rect 3936 4440 5356 4468
rect 3936 4428 3942 4440
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5534 4428 5540 4480
rect 5592 4428 5598 4480
rect 5994 4428 6000 4480
rect 6052 4428 6058 4480
rect 8110 4428 8116 4480
rect 8168 4428 8174 4480
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8294 4468 8300 4480
rect 8251 4440 8300 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8404 4468 8432 4508
rect 8478 4496 8484 4548
rect 8536 4496 8542 4548
rect 9582 4496 9588 4548
rect 9640 4508 9674 4548
rect 9769 4539 9827 4545
rect 9640 4496 9646 4508
rect 9769 4505 9781 4539
rect 9815 4536 9827 4539
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9815 4508 10149 4536
rect 9815 4505 9827 4508
rect 9769 4499 9827 4505
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10137 4499 10195 4505
rect 9858 4468 9864 4480
rect 8404 4440 9864 4468
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4468 11391 4471
rect 11606 4468 11612 4480
rect 11379 4440 11612 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 1104 4378 13984 4400
rect 1104 4326 4918 4378
rect 4970 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 5238 4378
rect 5290 4326 10918 4378
rect 10970 4326 10982 4378
rect 11034 4326 11046 4378
rect 11098 4326 11110 4378
rect 11162 4326 11174 4378
rect 11226 4326 11238 4378
rect 11290 4326 13984 4378
rect 1104 4304 13984 4326
rect 3418 4224 3424 4276
rect 3476 4224 3482 4276
rect 3878 4264 3884 4276
rect 3712 4236 3884 4264
rect 3712 4205 3740 4236
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5442 4264 5448 4276
rect 4488 4236 5448 4264
rect 4488 4224 4494 4236
rect 3053 4199 3111 4205
rect 3053 4165 3065 4199
rect 3099 4196 3111 4199
rect 3697 4199 3755 4205
rect 3697 4196 3709 4199
rect 3099 4168 3709 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 3697 4165 3709 4168
rect 3743 4196 3755 4199
rect 4341 4199 4399 4205
rect 4341 4196 4353 4199
rect 3743 4168 4353 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 4341 4165 4353 4168
rect 4387 4165 4399 4199
rect 4341 4159 4399 4165
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 2958 4128 2964 4140
rect 2915 4100 2964 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3142 4088 3148 4140
rect 3200 4088 3206 4140
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3252 3924 3280 4091
rect 3510 4088 3516 4140
rect 3568 4088 3574 4140
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 3970 4128 3976 4140
rect 3927 4100 3976 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 3804 3992 3832 4091
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4172 4060 4200 4091
rect 4430 4088 4436 4140
rect 4488 4088 4494 4140
rect 4540 4137 4568 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 6730 4224 6736 4276
rect 6788 4224 6794 4276
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8478 4264 8484 4276
rect 8435 4236 8484 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8478 4224 8484 4236
rect 8536 4264 8542 4276
rect 8536 4236 9536 4264
rect 8536 4224 8542 4236
rect 5258 4196 5264 4208
rect 4816 4168 5264 4196
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4816 4069 4844 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5057 4131 5115 4137
rect 5057 4128 5069 4131
rect 4948 4100 5069 4128
rect 4948 4088 4954 4100
rect 5057 4097 5069 4100
rect 5103 4097 5115 4131
rect 5552 4128 5580 4224
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 5552 4100 6561 4128
rect 5057 4091 5115 4097
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 4801 4063 4859 4069
rect 4172 4032 4384 4060
rect 4356 3992 4384 4032
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 6365 4063 6423 4069
rect 6365 4029 6377 4063
rect 6411 4060 6423 4063
rect 6748 4060 6776 4224
rect 9508 4208 9536 4236
rect 9582 4224 9588 4276
rect 9640 4224 9646 4276
rect 10042 4264 10048 4276
rect 9692 4236 10048 4264
rect 8665 4199 8723 4205
rect 8665 4196 8677 4199
rect 8312 4168 8677 4196
rect 8312 4140 8340 4168
rect 8665 4165 8677 4168
rect 8711 4165 8723 4199
rect 8665 4159 8723 4165
rect 9490 4156 9496 4208
rect 9548 4156 9554 4208
rect 9692 4196 9720 4236
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 11057 4267 11115 4273
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11330 4264 11336 4276
rect 11103 4236 11336 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 9600 4168 9720 4196
rect 9876 4168 10180 4196
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8110 4128 8116 4140
rect 6972 4100 8116 4128
rect 6972 4088 6978 4100
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8294 4128 8300 4140
rect 8251 4100 8300 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9401 4131 9459 4137
rect 8895 4100 9168 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 6411 4032 6776 4060
rect 6411 4029 6423 4032
rect 6365 4023 6423 4029
rect 6181 3995 6239 4001
rect 3804 3964 4292 3992
rect 4356 3964 4844 3992
rect 3970 3924 3976 3936
rect 3252 3896 3976 3924
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4062 3884 4068 3936
rect 4120 3884 4126 3936
rect 4264 3924 4292 3964
rect 4338 3924 4344 3936
rect 4264 3896 4344 3924
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 4706 3884 4712 3936
rect 4764 3884 4770 3936
rect 4816 3924 4844 3964
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 8496 3992 8524 4091
rect 9140 4069 9168 4100
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9600 4128 9628 4168
rect 9447 4100 9628 4128
rect 9677 4131 9735 4137
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 9876 4128 9904 4168
rect 9950 4137 9956 4140
rect 9723 4100 9904 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 9944 4091 9956 4137
rect 10008 4128 10014 4140
rect 10152 4128 10180 4168
rect 11532 4168 12204 4196
rect 11532 4137 11560 4168
rect 12176 4140 12204 4168
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10008 4100 10044 4128
rect 10152 4100 11529 4128
rect 9950 4088 9956 4091
rect 10008 4088 10014 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 11773 4131 11831 4137
rect 11773 4128 11785 4131
rect 11664 4100 11785 4128
rect 11664 4088 11670 4100
rect 11773 4097 11785 4100
rect 11819 4097 11831 4131
rect 11773 4091 11831 4097
rect 12158 4088 12164 4140
rect 12216 4088 12222 4140
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4060 9183 4063
rect 9214 4060 9220 4072
rect 9171 4032 9220 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 8662 3992 8668 4004
rect 6227 3964 8156 3992
rect 8496 3964 8668 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6196 3924 6224 3955
rect 4816 3896 6224 3924
rect 6733 3927 6791 3933
rect 6733 3893 6745 3927
rect 6779 3924 6791 3927
rect 7098 3924 7104 3936
rect 6779 3896 7104 3924
rect 6779 3893 6791 3896
rect 6733 3887 6791 3893
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 7708 3896 8033 3924
rect 7708 3884 7714 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8128 3924 8156 3964
rect 8662 3952 8668 3964
rect 8720 3992 8726 4004
rect 8720 3964 9168 3992
rect 8720 3952 8726 3964
rect 9140 3936 9168 3964
rect 8478 3924 8484 3936
rect 8128 3896 8484 3924
rect 8021 3887 8079 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 9030 3884 9036 3936
rect 9088 3884 9094 3936
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 9180 3896 9229 3924
rect 9180 3884 9186 3896
rect 9217 3893 9229 3896
rect 9263 3893 9275 3927
rect 9217 3887 9275 3893
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 11756 3896 12909 3924
rect 11756 3884 11762 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 1104 3834 13984 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13984 3834
rect 1104 3760 13984 3782
rect 3786 3720 3792 3732
rect 1964 3692 3792 3720
rect 1964 3525 1992 3692
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4062 3680 4068 3732
rect 4120 3680 4126 3732
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 4890 3720 4896 3732
rect 4479 3692 4896 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5537 3723 5595 3729
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5810 3720 5816 3732
rect 5583 3692 5816 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 10134 3680 10140 3732
rect 10192 3680 10198 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 13228 3692 13461 3720
rect 13228 3680 13234 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 3510 3612 3516 3664
rect 3568 3652 3574 3664
rect 3605 3655 3663 3661
rect 3605 3652 3617 3655
rect 3568 3624 3617 3652
rect 3568 3612 3574 3624
rect 3605 3621 3617 3624
rect 3651 3652 3663 3655
rect 3651 3624 3924 3652
rect 3651 3621 3663 3624
rect 3605 3615 3663 3621
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2314 3516 2320 3528
rect 2271 3488 2320 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2492 3451 2550 3457
rect 2492 3417 2504 3451
rect 2538 3448 2550 3451
rect 3694 3448 3700 3460
rect 2538 3420 3700 3448
rect 2538 3417 2550 3420
rect 2492 3411 2550 3417
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 3896 3448 3924 3624
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4080 3516 4108 3680
rect 4246 3612 4252 3664
rect 4304 3652 4310 3664
rect 5350 3652 5356 3664
rect 4304 3624 5120 3652
rect 4304 3612 4310 3624
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3584 4215 3587
rect 4614 3584 4620 3596
rect 4203 3556 4620 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 4614 3544 4620 3556
rect 4672 3584 4678 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4672 3556 4905 3584
rect 4672 3544 4678 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 4019 3488 4108 3516
rect 4249 3519 4307 3525
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4295 3488 4537 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 3896 3420 4752 3448
rect 4724 3392 4752 3420
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3380 2191 3383
rect 2314 3380 2320 3392
rect 2179 3352 2320 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 4706 3340 4712 3392
rect 4764 3340 4770 3392
rect 5000 3380 5028 3479
rect 5092 3448 5120 3624
rect 5184 3624 5356 3652
rect 5184 3525 5212 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 7009 3587 7067 3593
rect 5316 3556 5580 3584
rect 5316 3544 5322 3556
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5442 3516 5448 3528
rect 5399 3488 5448 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5552 3516 5580 3556
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7377 3587 7435 3593
rect 7377 3584 7389 3587
rect 7055 3556 7389 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7377 3553 7389 3556
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 5626 3516 5632 3528
rect 5552 3488 5632 3516
rect 5626 3476 5632 3488
rect 5684 3516 5690 3528
rect 6270 3516 6276 3528
rect 5684 3488 6276 3516
rect 5684 3476 5690 3488
rect 6270 3476 6276 3488
rect 6328 3516 6334 3528
rect 7024 3516 7052 3547
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 9950 3584 9956 3596
rect 8536 3556 9956 3584
rect 8536 3544 8542 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 6328 3488 7052 3516
rect 6328 3476 6334 3488
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7650 3525 7656 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7156 3488 7297 3516
rect 7156 3476 7162 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7644 3516 7656 3525
rect 7611 3488 7656 3516
rect 7285 3479 7343 3485
rect 7644 3479 7656 3488
rect 7650 3476 7656 3479
rect 7708 3476 7714 3528
rect 10152 3516 10180 3680
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10152 3488 10425 3516
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 12158 3516 12164 3528
rect 12115 3488 12164 3516
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 5261 3451 5319 3457
rect 5261 3448 5273 3451
rect 5092 3420 5273 3448
rect 5261 3417 5273 3420
rect 5307 3417 5319 3451
rect 5261 3411 5319 3417
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 6742 3451 6800 3457
rect 6742 3448 6754 3451
rect 6604 3420 6754 3448
rect 6604 3408 6610 3420
rect 6742 3417 6754 3420
rect 6788 3417 6800 3451
rect 6742 3411 6800 3417
rect 12336 3451 12394 3457
rect 12336 3417 12348 3451
rect 12382 3448 12394 3451
rect 13446 3448 13452 3460
rect 12382 3420 13452 3448
rect 12382 3417 12394 3420
rect 12336 3411 12394 3417
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 5626 3380 5632 3392
rect 5000 3352 5632 3380
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 7098 3340 7104 3392
rect 7156 3340 7162 3392
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 1104 3290 13984 3312
rect 1104 3238 4918 3290
rect 4970 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 5238 3290
rect 5290 3238 10918 3290
rect 10970 3238 10982 3290
rect 11034 3238 11046 3290
rect 11098 3238 11110 3290
rect 11162 3238 11174 3290
rect 11226 3238 11238 3290
rect 11290 3238 13984 3290
rect 1104 3216 13984 3238
rect 3694 3136 3700 3188
rect 3752 3136 3758 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5442 3176 5448 3188
rect 4856 3148 5448 3176
rect 4856 3136 4862 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6052 3148 6408 3176
rect 6052 3136 6058 3148
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2481 3043 2539 3049
rect 2481 3040 2493 3043
rect 2372 3012 2493 3040
rect 2372 3000 2378 3012
rect 2481 3009 2493 3012
rect 2527 3009 2539 3043
rect 2481 3003 2539 3009
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3844 3012 3893 3040
rect 3844 3000 3850 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 5925 3043 5983 3049
rect 5925 3009 5937 3043
rect 5971 3040 5983 3043
rect 6181 3043 6239 3049
rect 5971 3012 6132 3040
rect 5971 3009 5983 3012
rect 5925 3003 5983 3009
rect 6104 2972 6132 3012
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 6270 3040 6276 3052
rect 6227 3012 6276 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6380 3049 6408 3148
rect 6546 3136 6552 3188
rect 6604 3136 6610 3188
rect 7098 3136 7104 3188
rect 7156 3136 7162 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 9030 3136 9036 3188
rect 9088 3136 9094 3188
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 7116 2972 7144 3136
rect 7392 3040 7420 3136
rect 9048 3108 9076 3136
rect 8404 3080 9076 3108
rect 8404 3049 8432 3080
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7392 3012 8217 3040
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3009 8447 3043
rect 8389 3003 8447 3009
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8628 3012 8677 3040
rect 8628 3000 8634 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 10054 3043 10112 3049
rect 10054 3040 10066 3043
rect 8895 3012 10066 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 10054 3009 10066 3012
rect 10100 3009 10112 3043
rect 10054 3003 10112 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 12158 3040 12164 3052
rect 10367 3012 12164 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 6104 2944 7144 2972
rect 8404 2944 8616 2972
rect 8404 2916 8432 2944
rect 8386 2864 8392 2916
rect 8444 2864 8450 2916
rect 8478 2864 8484 2916
rect 8536 2864 8542 2916
rect 8588 2913 8616 2944
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3016 2808 3617 2836
rect 3016 2796 3022 2808
rect 3605 2805 3617 2808
rect 3651 2836 3663 2839
rect 5534 2836 5540 2848
rect 3651 2808 5540 2836
rect 3651 2805 3663 2808
rect 3605 2799 3663 2805
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 8941 2839 8999 2845
rect 8941 2805 8953 2839
rect 8987 2836 8999 2839
rect 9214 2836 9220 2848
rect 8987 2808 9220 2836
rect 8987 2805 8999 2808
rect 8941 2799 8999 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 1104 2746 13984 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13984 2746
rect 1104 2672 13984 2694
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8536 2604 9137 2632
rect 8536 2592 8542 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 9490 2592 9496 2644
rect 9548 2632 9554 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 9548 2604 9597 2632
rect 9548 2592 9554 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 13446 2592 13452 2644
rect 13504 2592 13510 2644
rect 8754 2524 8760 2576
rect 8812 2524 8818 2576
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 9769 2567 9827 2573
rect 9769 2564 9781 2567
rect 9364 2536 9781 2564
rect 9364 2524 9370 2536
rect 9769 2533 9781 2536
rect 9815 2533 9827 2567
rect 9769 2527 9827 2533
rect 2866 2496 2872 2508
rect 1596 2468 2872 2496
rect 1596 2437 1624 2468
rect 2866 2456 2872 2468
rect 2924 2456 2930 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5684 2468 8432 2496
rect 5684 2456 5690 2468
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 1728 2400 2421 2428
rect 1728 2388 1734 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 3602 2388 3608 2440
rect 3660 2388 3666 2440
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 8404 2437 8432 2468
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5592 2400 6009 2428
rect 5592 2388 5598 2400
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 5997 2391 6055 2397
rect 6886 2400 7205 2428
rect 5442 2320 5448 2372
rect 5500 2360 5506 2372
rect 6886 2360 6914 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8772 2428 8800 2524
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 8772 2400 9413 2428
rect 8389 2391 8447 2397
rect 9401 2397 9413 2400
rect 9447 2428 9459 2431
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9447 2400 9505 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10652 2400 10793 2428
rect 10652 2388 10658 2400
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11756 2400 11989 2428
rect 11756 2388 11762 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13354 2428 13360 2440
rect 13219 2400 13360 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 14090 2428 14096 2440
rect 13679 2400 14096 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 5500 2332 6914 2360
rect 5500 2320 5506 2332
rect 9122 2320 9128 2372
rect 9180 2320 9186 2372
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 9272 2332 9321 2360
rect 9272 2320 9278 2332
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9309 2323 9367 2329
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 992 2264 1409 2292
rect 992 2252 998 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 2222 2252 2228 2304
rect 2280 2252 2286 2304
rect 3418 2252 3424 2304
rect 3476 2252 3482 2304
rect 4614 2252 4620 2304
rect 4672 2252 4678 2304
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 7006 2252 7012 2304
rect 7064 2252 7070 2304
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 10594 2252 10600 2304
rect 10652 2252 10658 2304
rect 11790 2252 11796 2304
rect 11848 2252 11854 2304
rect 12986 2252 12992 2304
rect 13044 2252 13050 2304
rect 1104 2202 13984 2224
rect 1104 2150 4918 2202
rect 4970 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 5238 2202
rect 5290 2150 10918 2202
rect 10970 2150 10982 2202
rect 11034 2150 11046 2202
rect 11098 2150 11110 2202
rect 11162 2150 11174 2202
rect 11226 2150 11238 2202
rect 11290 2150 13984 2202
rect 1104 2128 13984 2150
<< via1 >>
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 940 14560 992 14612
rect 2320 14560 2372 14612
rect 3056 14603 3108 14612
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 3976 14560 4028 14612
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 6000 14560 6052 14612
rect 7012 14560 7064 14612
rect 7840 14560 7892 14612
rect 9036 14560 9088 14612
rect 3516 14492 3568 14544
rect 5448 14492 5500 14544
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 2780 14356 2832 14408
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 3700 14288 3752 14340
rect 5356 14356 5408 14408
rect 7748 14356 7800 14408
rect 11060 14356 11112 14408
rect 12072 14356 12124 14408
rect 13084 14356 13136 14408
rect 5632 14220 5684 14272
rect 6920 14220 6972 14272
rect 8576 14220 8628 14272
rect 11336 14263 11388 14272
rect 11336 14229 11345 14263
rect 11345 14229 11379 14263
rect 11379 14229 11388 14263
rect 11336 14220 11388 14229
rect 11888 14220 11940 14272
rect 4918 14118 4970 14170
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 5238 14118 5290 14170
rect 10918 14118 10970 14170
rect 10982 14118 11034 14170
rect 11046 14118 11098 14170
rect 11110 14118 11162 14170
rect 11174 14118 11226 14170
rect 11238 14118 11290 14170
rect 6920 14016 6972 14068
rect 2872 13880 2924 13932
rect 2964 13880 3016 13932
rect 3516 13880 3568 13932
rect 3792 13880 3844 13932
rect 4068 13880 4120 13932
rect 4436 13948 4488 14000
rect 5356 13948 5408 14000
rect 4528 13880 4580 13932
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 7104 13991 7156 14000
rect 7104 13957 7113 13991
rect 7113 13957 7147 13991
rect 7147 13957 7156 13991
rect 7104 13948 7156 13957
rect 7748 13948 7800 14000
rect 7196 13880 7248 13932
rect 8668 13880 8720 13932
rect 9772 13880 9824 13932
rect 10140 13880 10192 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 11520 13880 11572 13932
rect 6644 13812 6696 13864
rect 6828 13812 6880 13864
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 4804 13744 4856 13796
rect 9680 13812 9732 13864
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 6184 13676 6236 13728
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 3976 13472 4028 13524
rect 4068 13472 4120 13524
rect 5632 13472 5684 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 6368 13472 6420 13524
rect 6736 13472 6788 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 3056 13404 3108 13456
rect 3700 13404 3752 13456
rect 5448 13404 5500 13456
rect 8668 13472 8720 13524
rect 2688 13268 2740 13320
rect 3332 13268 3384 13320
rect 6184 13336 6236 13388
rect 5724 13268 5776 13320
rect 6736 13336 6788 13388
rect 7196 13311 7248 13320
rect 7196 13277 7205 13311
rect 7205 13277 7239 13311
rect 7239 13277 7248 13311
rect 7196 13268 7248 13277
rect 9680 13268 9732 13320
rect 12072 13268 12124 13320
rect 2136 13200 2188 13252
rect 2872 13132 2924 13184
rect 2964 13132 3016 13184
rect 5356 13243 5408 13252
rect 5356 13209 5365 13243
rect 5365 13209 5399 13243
rect 5399 13209 5408 13243
rect 5356 13200 5408 13209
rect 6368 13200 6420 13252
rect 3884 13132 3936 13184
rect 6460 13132 6512 13184
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 10692 13243 10744 13252
rect 10692 13209 10726 13243
rect 10726 13209 10744 13243
rect 10692 13200 10744 13209
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 9220 13132 9272 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 4918 13030 4970 13082
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 5238 13030 5290 13082
rect 10918 13030 10970 13082
rect 10982 13030 11034 13082
rect 11046 13030 11098 13082
rect 11110 13030 11162 13082
rect 11174 13030 11226 13082
rect 11238 13030 11290 13082
rect 2136 12971 2188 12980
rect 2136 12937 2145 12971
rect 2145 12937 2179 12971
rect 2179 12937 2188 12971
rect 2136 12928 2188 12937
rect 2872 12928 2924 12980
rect 3884 12928 3936 12980
rect 4528 12928 4580 12980
rect 4804 12928 4856 12980
rect 2320 12835 2372 12844
rect 2320 12801 2329 12835
rect 2329 12801 2363 12835
rect 2363 12801 2372 12835
rect 2320 12792 2372 12801
rect 3332 12792 3384 12844
rect 5816 12928 5868 12980
rect 7196 12928 7248 12980
rect 7748 12928 7800 12980
rect 9772 12928 9824 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 11796 12928 11848 12980
rect 5264 12903 5316 12912
rect 5264 12869 5273 12903
rect 5273 12869 5307 12903
rect 5307 12869 5316 12903
rect 5264 12860 5316 12869
rect 8944 12860 8996 12912
rect 10600 12860 10652 12912
rect 2688 12724 2740 12776
rect 6276 12724 6328 12776
rect 9496 12792 9548 12844
rect 8668 12724 8720 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 3976 12588 4028 12640
rect 5264 12656 5316 12708
rect 10416 12724 10468 12776
rect 11612 12792 11664 12844
rect 5356 12588 5408 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 9772 12588 9824 12640
rect 11336 12656 11388 12708
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 12440 12656 12492 12708
rect 12532 12656 12584 12708
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 3700 12316 3752 12368
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 4712 12316 4764 12368
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 6000 12427 6052 12436
rect 6000 12393 6021 12427
rect 6021 12393 6052 12427
rect 6000 12384 6052 12393
rect 6092 12384 6144 12436
rect 6736 12427 6788 12436
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 9864 12384 9916 12436
rect 9956 12384 10008 12436
rect 8668 12316 8720 12368
rect 2964 12248 3016 12257
rect 4804 12248 4856 12300
rect 2504 12155 2556 12164
rect 2504 12121 2513 12155
rect 2513 12121 2547 12155
rect 2547 12121 2556 12155
rect 2504 12112 2556 12121
rect 1676 12044 1728 12096
rect 2596 12044 2648 12096
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3240 12180 3292 12232
rect 4252 12112 4304 12164
rect 5540 12180 5592 12232
rect 5816 12180 5868 12232
rect 5908 12180 5960 12232
rect 6184 12155 6236 12164
rect 6184 12121 6193 12155
rect 6193 12121 6227 12155
rect 6227 12121 6236 12155
rect 6184 12112 6236 12121
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9680 12180 9732 12232
rect 9956 12223 10008 12232
rect 9956 12189 9960 12223
rect 9960 12189 9994 12223
rect 9994 12189 10008 12223
rect 9956 12180 10008 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 10968 12248 11020 12300
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 7104 12112 7156 12164
rect 3056 12044 3108 12096
rect 3332 12044 3384 12096
rect 3516 12044 3568 12096
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 5356 12044 5408 12096
rect 5724 12044 5776 12096
rect 9864 12112 9916 12164
rect 10048 12155 10100 12164
rect 10048 12121 10057 12155
rect 10057 12121 10091 12155
rect 10091 12121 10100 12155
rect 10048 12112 10100 12121
rect 10600 12112 10652 12164
rect 11244 12316 11296 12368
rect 11796 12316 11848 12368
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 11704 12248 11756 12300
rect 11336 12180 11388 12232
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 11244 12044 11296 12096
rect 11796 12044 11848 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12072 12044 12124 12096
rect 12256 12112 12308 12164
rect 12624 12044 12676 12096
rect 4918 11942 4970 11994
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 5238 11942 5290 11994
rect 10918 11942 10970 11994
rect 10982 11942 11034 11994
rect 11046 11942 11098 11994
rect 11110 11942 11162 11994
rect 11174 11942 11226 11994
rect 11238 11942 11290 11994
rect 2504 11840 2556 11892
rect 2688 11772 2740 11824
rect 3240 11772 3292 11824
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 4436 11840 4488 11892
rect 1768 11747 1820 11756
rect 1768 11713 1802 11747
rect 1802 11713 1820 11747
rect 1768 11704 1820 11713
rect 2872 11636 2924 11688
rect 3332 11636 3384 11688
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 4436 11704 4488 11756
rect 4896 11772 4948 11824
rect 4988 11815 5040 11824
rect 4988 11781 4997 11815
rect 4997 11781 5031 11815
rect 5031 11781 5040 11815
rect 4988 11772 5040 11781
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 5356 11840 5408 11892
rect 3608 11636 3660 11645
rect 4252 11636 4304 11688
rect 4712 11636 4764 11688
rect 4804 11636 4856 11688
rect 5080 11636 5132 11688
rect 6000 11772 6052 11824
rect 10324 11840 10376 11892
rect 10692 11840 10744 11892
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 10876 11840 10928 11892
rect 11336 11840 11388 11892
rect 11612 11883 11664 11892
rect 11612 11849 11621 11883
rect 11621 11849 11655 11883
rect 11655 11849 11664 11883
rect 11612 11840 11664 11849
rect 11796 11840 11848 11892
rect 11980 11840 12032 11892
rect 12164 11840 12216 11892
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 6092 11636 6144 11688
rect 2780 11500 2832 11552
rect 4252 11500 4304 11552
rect 5816 11500 5868 11552
rect 6276 11568 6328 11620
rect 9404 11772 9456 11824
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 9772 11772 9824 11824
rect 9588 11704 9640 11756
rect 10048 11704 10100 11756
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 6552 11636 6604 11688
rect 6828 11636 6880 11688
rect 7288 11679 7340 11688
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7472 11636 7524 11688
rect 9312 11636 9364 11688
rect 6920 11568 6972 11620
rect 7840 11611 7892 11620
rect 7840 11577 7849 11611
rect 7849 11577 7883 11611
rect 7883 11577 7892 11611
rect 7840 11568 7892 11577
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 12256 11815 12308 11824
rect 12256 11781 12265 11815
rect 12265 11781 12299 11815
rect 12299 11781 12308 11815
rect 12256 11772 12308 11781
rect 12440 11840 12492 11892
rect 12624 11772 12676 11824
rect 11244 11568 11296 11620
rect 11336 11568 11388 11620
rect 11612 11568 11664 11620
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 6460 11500 6512 11552
rect 7012 11500 7064 11552
rect 8668 11500 8720 11552
rect 9220 11500 9272 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 9956 11500 10008 11552
rect 10416 11500 10468 11552
rect 10968 11500 11020 11552
rect 11060 11500 11112 11552
rect 12164 11500 12216 11552
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 1768 11296 1820 11348
rect 2320 11296 2372 11348
rect 2596 11296 2648 11348
rect 1676 11160 1728 11212
rect 3332 11228 3384 11280
rect 3056 11160 3108 11212
rect 4344 11296 4396 11348
rect 3976 11228 4028 11280
rect 4896 11228 4948 11280
rect 4344 11092 4396 11144
rect 4712 11092 4764 11144
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5172 11296 5224 11348
rect 6368 11296 6420 11348
rect 6552 11296 6604 11348
rect 6920 11296 6972 11348
rect 7104 11339 7156 11348
rect 7104 11305 7113 11339
rect 7113 11305 7147 11339
rect 7147 11305 7156 11339
rect 7104 11296 7156 11305
rect 7748 11296 7800 11348
rect 5632 11228 5684 11280
rect 3240 11024 3292 11076
rect 2872 10956 2924 11008
rect 4068 10956 4120 11008
rect 4160 10999 4212 11008
rect 4160 10965 4169 10999
rect 4169 10965 4203 10999
rect 4203 10965 4212 10999
rect 4160 10956 4212 10965
rect 4712 10956 4764 11008
rect 4804 10956 4856 11008
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 5908 11160 5960 11212
rect 6000 11160 6052 11212
rect 6184 11160 6236 11212
rect 5632 11135 5684 11144
rect 5632 11101 5641 11135
rect 5641 11101 5675 11135
rect 5675 11101 5684 11135
rect 5632 11092 5684 11101
rect 7472 11271 7524 11280
rect 7472 11237 7481 11271
rect 7481 11237 7515 11271
rect 7515 11237 7524 11271
rect 7472 11228 7524 11237
rect 7656 11228 7708 11280
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6736 11092 6788 11144
rect 7932 11092 7984 11144
rect 8300 11092 8352 11144
rect 8944 11296 8996 11348
rect 10600 11296 10652 11348
rect 8668 11271 8720 11280
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 11244 11228 11296 11280
rect 11428 11296 11480 11348
rect 11612 11228 11664 11280
rect 11336 11160 11388 11212
rect 11980 11228 12032 11280
rect 9220 11092 9272 11144
rect 6276 11024 6328 11076
rect 7288 11024 7340 11076
rect 7380 11024 7432 11076
rect 8392 11067 8444 11076
rect 8392 11033 8401 11067
rect 8401 11033 8435 11067
rect 8435 11033 8444 11067
rect 8392 11024 8444 11033
rect 10324 11024 10376 11076
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 11428 11092 11480 11144
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 6736 10956 6788 11008
rect 7932 10956 7984 11008
rect 8576 10956 8628 11008
rect 10968 10956 11020 11008
rect 11612 10956 11664 11008
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 12072 10956 12124 11008
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 12716 10956 12768 11008
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 4918 10854 4970 10906
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 5238 10854 5290 10906
rect 10918 10854 10970 10906
rect 10982 10854 11034 10906
rect 11046 10854 11098 10906
rect 11110 10854 11162 10906
rect 11174 10854 11226 10906
rect 11238 10854 11290 10906
rect 3608 10795 3660 10804
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4068 10795 4120 10804
rect 4068 10761 4077 10795
rect 4077 10761 4111 10795
rect 4111 10761 4120 10795
rect 4068 10752 4120 10761
rect 4528 10752 4580 10804
rect 4344 10684 4396 10736
rect 4160 10616 4212 10668
rect 4620 10616 4672 10668
rect 4896 10616 4948 10668
rect 5356 10752 5408 10804
rect 6368 10752 6420 10804
rect 7380 10752 7432 10804
rect 7472 10752 7524 10804
rect 8024 10752 8076 10804
rect 9772 10752 9824 10804
rect 6644 10684 6696 10736
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 6000 10616 6052 10668
rect 6552 10616 6604 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7656 10616 7708 10668
rect 8300 10616 8352 10668
rect 4804 10480 4856 10532
rect 4620 10412 4672 10464
rect 6644 10548 6696 10600
rect 7288 10548 7340 10600
rect 8576 10616 8628 10668
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9404 10616 9456 10668
rect 6368 10480 6420 10532
rect 10048 10684 10100 10736
rect 11152 10752 11204 10804
rect 12072 10752 12124 10804
rect 12164 10752 12216 10804
rect 10600 10616 10652 10668
rect 10784 10616 10836 10668
rect 11060 10616 11112 10668
rect 11244 10684 11296 10736
rect 12716 10684 12768 10736
rect 10048 10548 10100 10600
rect 11612 10548 11664 10600
rect 12992 10616 13044 10668
rect 9588 10523 9640 10532
rect 9588 10489 9597 10523
rect 9597 10489 9631 10523
rect 9631 10489 9640 10523
rect 9588 10480 9640 10489
rect 9680 10480 9732 10532
rect 10784 10523 10836 10532
rect 10784 10489 10793 10523
rect 10793 10489 10827 10523
rect 10827 10489 10836 10523
rect 10784 10480 10836 10489
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 6828 10412 6880 10464
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 7748 10412 7800 10421
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 10140 10412 10192 10464
rect 10324 10412 10376 10464
rect 12072 10480 12124 10532
rect 13176 10548 13228 10600
rect 11152 10412 11204 10464
rect 11428 10412 11480 10464
rect 12164 10412 12216 10464
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 4712 10208 4764 10260
rect 5816 10208 5868 10260
rect 4896 10140 4948 10192
rect 6552 10140 6604 10192
rect 6828 10208 6880 10260
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7196 10208 7248 10260
rect 7840 10251 7892 10260
rect 7840 10217 7849 10251
rect 7849 10217 7883 10251
rect 7883 10217 7892 10251
rect 7840 10208 7892 10217
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 9036 10208 9088 10260
rect 6736 10140 6788 10192
rect 11704 10208 11756 10260
rect 12532 10140 12584 10192
rect 6644 10072 6696 10124
rect 3976 10004 4028 10056
rect 6460 10004 6512 10056
rect 6828 10004 6880 10056
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7196 10115 7248 10124
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 7656 10072 7708 10124
rect 7380 10004 7432 10056
rect 7472 10004 7524 10056
rect 11704 10072 11756 10124
rect 11796 10072 11848 10124
rect 8576 10047 8628 10056
rect 7840 9936 7892 9988
rect 4344 9868 4396 9920
rect 6368 9868 6420 9920
rect 7288 9868 7340 9920
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8392 9936 8444 9988
rect 10692 10004 10744 10056
rect 11060 10004 11112 10056
rect 12164 10004 12216 10056
rect 12992 10004 13044 10056
rect 10048 9979 10100 9988
rect 10048 9945 10066 9979
rect 10066 9945 10100 9979
rect 10048 9936 10100 9945
rect 8484 9868 8536 9920
rect 9036 9868 9088 9920
rect 9128 9868 9180 9920
rect 12624 9936 12676 9988
rect 10692 9868 10744 9920
rect 11244 9868 11296 9920
rect 12256 9868 12308 9920
rect 4918 9766 4970 9818
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 5238 9766 5290 9818
rect 10918 9766 10970 9818
rect 10982 9766 11034 9818
rect 11046 9766 11098 9818
rect 11110 9766 11162 9818
rect 11174 9766 11226 9818
rect 11238 9766 11290 9818
rect 4804 9664 4856 9716
rect 2780 9596 2832 9648
rect 4344 9596 4396 9648
rect 3424 9528 3476 9580
rect 4160 9528 4212 9580
rect 5908 9596 5960 9648
rect 6736 9596 6788 9648
rect 7840 9664 7892 9716
rect 9128 9664 9180 9716
rect 9404 9664 9456 9716
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 10140 9664 10192 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 10508 9664 10560 9716
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 2964 9460 3016 9512
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3516 9460 3568 9512
rect 3884 9460 3936 9512
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 6920 9460 6972 9512
rect 3240 9392 3292 9444
rect 3976 9324 4028 9376
rect 7104 9392 7156 9444
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 11704 9664 11756 9716
rect 11796 9664 11848 9716
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 9128 9392 9180 9444
rect 9680 9392 9732 9444
rect 9772 9392 9824 9444
rect 10692 9460 10744 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11244 9596 11296 9648
rect 11428 9528 11480 9580
rect 11796 9528 11848 9580
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 6276 9324 6328 9376
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 7380 9324 7432 9376
rect 8944 9324 8996 9376
rect 13360 9392 13412 9444
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 10968 9324 11020 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 1584 9120 1636 9172
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 3056 9120 3108 9172
rect 3240 9120 3292 9172
rect 4252 9120 4304 9172
rect 4620 9120 4672 9172
rect 3332 9052 3384 9104
rect 4712 9052 4764 9104
rect 1676 8916 1728 8968
rect 2780 8916 2832 8968
rect 1952 8848 2004 8900
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3332 8916 3384 8968
rect 3884 8916 3936 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 5816 9052 5868 9104
rect 5448 8984 5500 9036
rect 7196 9120 7248 9172
rect 7472 9120 7524 9172
rect 9404 9120 9456 9172
rect 9588 9120 9640 9172
rect 2872 8780 2924 8832
rect 3240 8780 3292 8832
rect 3424 8780 3476 8832
rect 4528 8848 4580 8900
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5632 8916 5684 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6368 8916 6420 8968
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 3884 8780 3936 8832
rect 6276 8780 6328 8832
rect 6552 8848 6604 8900
rect 8760 8916 8812 8968
rect 6920 8848 6972 8900
rect 9772 8984 9824 9036
rect 10416 9120 10468 9172
rect 10876 9120 10928 9172
rect 11060 9052 11112 9104
rect 12716 9120 12768 9172
rect 10600 8984 10652 9036
rect 9128 8916 9180 8968
rect 9864 8916 9916 8968
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 10876 8984 10928 9036
rect 11244 8984 11296 9036
rect 11336 8984 11388 9036
rect 9772 8848 9824 8900
rect 6644 8780 6696 8832
rect 7748 8780 7800 8832
rect 9680 8780 9732 8832
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 10508 8780 10560 8832
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11704 8984 11756 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 11980 8916 12032 8968
rect 12164 8848 12216 8900
rect 12532 8848 12584 8900
rect 12992 8780 13044 8832
rect 4918 8678 4970 8730
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 5238 8678 5290 8730
rect 10918 8678 10970 8730
rect 10982 8678 11034 8730
rect 11046 8678 11098 8730
rect 11110 8678 11162 8730
rect 11174 8678 11226 8730
rect 11238 8678 11290 8730
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 1584 8440 1636 8492
rect 3976 8576 4028 8628
rect 4252 8576 4304 8628
rect 5816 8576 5868 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 6460 8576 6512 8628
rect 6644 8576 6696 8628
rect 4528 8551 4580 8560
rect 4528 8517 4537 8551
rect 4537 8517 4571 8551
rect 4571 8517 4580 8551
rect 4528 8508 4580 8517
rect 6276 8508 6328 8560
rect 7564 8576 7616 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8760 8576 8812 8628
rect 11428 8576 11480 8628
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 2780 8440 2832 8492
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2872 8372 2924 8424
rect 2964 8304 3016 8356
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 6552 8440 6604 8492
rect 6920 8440 6972 8492
rect 5632 8372 5684 8424
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 7748 8440 7800 8492
rect 5908 8372 5960 8381
rect 5172 8304 5224 8356
rect 5356 8304 5408 8356
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 5080 8236 5132 8288
rect 5724 8236 5776 8288
rect 6828 8236 6880 8288
rect 7104 8236 7156 8288
rect 14096 8508 14148 8560
rect 9864 8440 9916 8492
rect 10508 8440 10560 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 11152 8440 11204 8492
rect 11612 8440 11664 8492
rect 9772 8372 9824 8424
rect 10876 8372 10928 8424
rect 10600 8304 10652 8356
rect 12256 8440 12308 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13360 8440 13412 8492
rect 9772 8236 9824 8288
rect 10232 8236 10284 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 4252 8032 4304 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5356 8032 5408 8084
rect 7196 8032 7248 8084
rect 7380 8032 7432 8084
rect 8392 8032 8444 8084
rect 3516 7964 3568 8016
rect 4068 7964 4120 8016
rect 4160 7964 4212 8016
rect 4804 7964 4856 8016
rect 5448 7964 5500 8016
rect 7748 7964 7800 8016
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 3424 7896 3476 7948
rect 4620 7896 4672 7948
rect 6184 7939 6236 7948
rect 6184 7905 6218 7939
rect 6218 7905 6236 7939
rect 6184 7896 6236 7905
rect 6368 7896 6420 7948
rect 6644 7896 6696 7948
rect 7380 7896 7432 7948
rect 4528 7828 4580 7880
rect 4712 7828 4764 7880
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 2964 7692 3016 7744
rect 3792 7760 3844 7812
rect 4252 7760 4304 7812
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 5448 7828 5500 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 5724 7871 5776 7880
rect 5724 7837 5740 7871
rect 5740 7837 5774 7871
rect 5774 7837 5776 7871
rect 5724 7828 5776 7837
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 7104 7828 7156 7880
rect 10048 8032 10100 8084
rect 10600 8032 10652 8084
rect 10784 8032 10836 8084
rect 8668 7896 8720 7948
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 3608 7692 3660 7744
rect 6000 7692 6052 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 8392 7692 8444 7744
rect 9772 7964 9824 8016
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10048 7692 10100 7744
rect 10876 7828 10928 7880
rect 4918 7590 4970 7642
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 5238 7590 5290 7642
rect 10918 7590 10970 7642
rect 10982 7590 11034 7642
rect 11046 7590 11098 7642
rect 11110 7590 11162 7642
rect 11174 7590 11226 7642
rect 11238 7590 11290 7642
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 6092 7488 6144 7540
rect 6736 7488 6788 7540
rect 7564 7531 7616 7540
rect 7564 7497 7573 7531
rect 7573 7497 7607 7531
rect 7607 7497 7616 7531
rect 7564 7488 7616 7497
rect 5356 7420 5408 7472
rect 5632 7352 5684 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6000 7395 6052 7404
rect 6000 7361 6006 7395
rect 6006 7361 6040 7395
rect 6040 7361 6052 7395
rect 7104 7420 7156 7472
rect 6000 7352 6052 7361
rect 6920 7352 6972 7404
rect 7288 7352 7340 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7472 7352 7524 7404
rect 7748 7352 7800 7404
rect 8668 7488 8720 7540
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 11520 7488 11572 7540
rect 8392 7463 8444 7472
rect 8392 7429 8401 7463
rect 8401 7429 8435 7463
rect 8435 7429 8444 7463
rect 8392 7420 8444 7429
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 6460 7327 6512 7336
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 6736 7284 6788 7336
rect 7656 7284 7708 7336
rect 5724 7216 5776 7268
rect 5816 7148 5868 7200
rect 6460 7148 6512 7200
rect 8576 7216 8628 7268
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 11428 7352 11480 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11888 7352 11940 7404
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 10048 7148 10100 7200
rect 10232 7148 10284 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 5908 6944 5960 6996
rect 7196 6944 7248 6996
rect 7748 6944 7800 6996
rect 9036 6987 9088 6996
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 3976 6808 4028 6860
rect 7288 6876 7340 6928
rect 7472 6808 7524 6860
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 9496 6944 9548 6996
rect 9864 6944 9916 6996
rect 8668 6876 8720 6928
rect 9956 6919 10008 6928
rect 9956 6885 9965 6919
rect 9965 6885 9999 6919
rect 9999 6885 10008 6919
rect 9956 6876 10008 6885
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 2964 6672 3016 6724
rect 4804 6740 4856 6792
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6920 6740 6972 6792
rect 7104 6740 7156 6792
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 4804 6604 4856 6656
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8024 6672 8076 6724
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9128 6672 9180 6724
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 10232 6808 10284 6860
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 9772 6715 9824 6724
rect 9772 6681 9781 6715
rect 9781 6681 9815 6715
rect 9815 6681 9824 6715
rect 9772 6672 9824 6681
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 8760 6604 8812 6656
rect 9312 6604 9364 6656
rect 10784 6740 10836 6792
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 11704 6740 11756 6792
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 13452 6740 13504 6792
rect 11336 6672 11388 6724
rect 10784 6604 10836 6656
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 4918 6502 4970 6554
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 5238 6502 5290 6554
rect 10918 6502 10970 6554
rect 10982 6502 11034 6554
rect 11046 6502 11098 6554
rect 11110 6502 11162 6554
rect 11174 6502 11226 6554
rect 11238 6502 11290 6554
rect 3056 6400 3108 6452
rect 3240 6400 3292 6452
rect 2964 6264 3016 6316
rect 3792 6400 3844 6452
rect 6276 6400 6328 6452
rect 8944 6400 8996 6452
rect 10048 6400 10100 6452
rect 6920 6332 6972 6384
rect 3608 6128 3660 6180
rect 1676 6060 1728 6112
rect 3976 6264 4028 6316
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 7472 6264 7524 6316
rect 8576 6375 8628 6384
rect 8576 6341 8585 6375
rect 8585 6341 8619 6375
rect 8619 6341 8628 6375
rect 8576 6332 8628 6341
rect 9036 6332 9088 6384
rect 9220 6332 9272 6384
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8300 6264 8352 6316
rect 8760 6264 8812 6316
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 11336 6400 11388 6452
rect 11428 6332 11480 6384
rect 4712 6196 4764 6248
rect 4528 6128 4580 6180
rect 8484 6196 8536 6248
rect 9036 6196 9088 6248
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10968 6264 11020 6316
rect 11336 6264 11388 6316
rect 7656 6171 7708 6180
rect 7656 6137 7665 6171
rect 7665 6137 7699 6171
rect 7699 6137 7708 6171
rect 7656 6128 7708 6137
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 4620 6060 4672 6112
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 8300 6060 8352 6112
rect 8484 6060 8536 6112
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 9312 6128 9364 6180
rect 13360 6196 13412 6248
rect 9404 6060 9456 6112
rect 9772 6060 9824 6112
rect 10968 6060 11020 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 2964 5856 3016 5908
rect 3332 5856 3384 5908
rect 3884 5856 3936 5908
rect 4068 5856 4120 5908
rect 7380 5856 7432 5908
rect 8392 5856 8444 5908
rect 10140 5856 10192 5908
rect 10968 5856 11020 5908
rect 2320 5652 2372 5704
rect 4436 5788 4488 5840
rect 7748 5788 7800 5840
rect 3608 5720 3660 5772
rect 3976 5720 4028 5772
rect 2964 5584 3016 5636
rect 3700 5584 3752 5636
rect 1768 5516 1820 5568
rect 3608 5559 3660 5568
rect 3608 5525 3617 5559
rect 3617 5525 3651 5559
rect 3651 5525 3660 5559
rect 3608 5516 3660 5525
rect 3884 5516 3936 5568
rect 9128 5788 9180 5840
rect 9588 5788 9640 5840
rect 7840 5652 7892 5704
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 9680 5720 9732 5772
rect 8484 5652 8536 5661
rect 6552 5584 6604 5636
rect 9036 5652 9088 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 4804 5516 4856 5568
rect 5632 5516 5684 5568
rect 9312 5516 9364 5568
rect 10048 5652 10100 5704
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 12072 5831 12124 5840
rect 12072 5797 12081 5831
rect 12081 5797 12115 5831
rect 12115 5797 12124 5831
rect 12072 5788 12124 5797
rect 12164 5652 12216 5704
rect 13360 5652 13412 5704
rect 13176 5627 13228 5636
rect 13176 5593 13194 5627
rect 13194 5593 13228 5627
rect 13176 5584 13228 5593
rect 4918 5414 4970 5466
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 5238 5414 5290 5466
rect 10918 5414 10970 5466
rect 10982 5414 11034 5466
rect 11046 5414 11098 5466
rect 11110 5414 11162 5466
rect 11174 5414 11226 5466
rect 11238 5414 11290 5466
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 3332 5312 3384 5364
rect 3884 5312 3936 5364
rect 4436 5355 4488 5364
rect 4436 5321 4445 5355
rect 4445 5321 4479 5355
rect 4479 5321 4488 5355
rect 4436 5312 4488 5321
rect 1768 5219 1820 5228
rect 1768 5185 1802 5219
rect 1802 5185 1820 5219
rect 1768 5176 1820 5185
rect 2320 5176 2372 5228
rect 4528 5244 4580 5296
rect 7380 5312 7432 5364
rect 6920 5244 6972 5296
rect 9036 5312 9088 5364
rect 9404 5312 9456 5364
rect 10784 5312 10836 5364
rect 11520 5312 11572 5364
rect 11796 5312 11848 5364
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 3976 5176 4028 5228
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 4712 5040 4764 5092
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 6460 5176 6512 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 8300 5244 8352 5296
rect 8392 5244 8444 5296
rect 7104 5176 7156 5228
rect 5724 5040 5776 5092
rect 6552 5040 6604 5092
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9128 5176 9180 5228
rect 9496 5244 9548 5296
rect 12348 5287 12400 5296
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 10232 5176 10284 5228
rect 11336 5176 11388 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12348 5253 12382 5287
rect 12382 5253 12400 5287
rect 12348 5244 12400 5253
rect 12164 5176 12216 5228
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 9312 4972 9364 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 6644 4768 6696 4820
rect 6736 4768 6788 4820
rect 9496 4768 9548 4820
rect 3424 4564 3476 4616
rect 4712 4564 4764 4616
rect 4804 4564 4856 4616
rect 4160 4496 4212 4548
rect 5540 4564 5592 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 9680 4700 9732 4752
rect 9956 4700 10008 4752
rect 7380 4632 7432 4684
rect 8392 4632 8444 4684
rect 9128 4632 9180 4684
rect 10692 4768 10744 4820
rect 11060 4768 11112 4820
rect 8576 4564 8628 4616
rect 9312 4564 9364 4616
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 3884 4428 3936 4480
rect 6736 4496 6788 4548
rect 5356 4428 5408 4480
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 8116 4428 8168 4480
rect 8300 4428 8352 4480
rect 8484 4539 8536 4548
rect 8484 4505 8493 4539
rect 8493 4505 8527 4539
rect 8527 4505 8536 4539
rect 8484 4496 8536 4505
rect 9588 4539 9640 4548
rect 9588 4505 9597 4539
rect 9597 4505 9631 4539
rect 9631 4505 9640 4539
rect 9588 4496 9640 4505
rect 9864 4428 9916 4480
rect 11612 4428 11664 4480
rect 4918 4326 4970 4378
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 5238 4326 5290 4378
rect 10918 4326 10970 4378
rect 10982 4326 11034 4378
rect 11046 4326 11098 4378
rect 11110 4326 11162 4378
rect 11174 4326 11226 4378
rect 11238 4326 11290 4378
rect 3424 4267 3476 4276
rect 3424 4233 3433 4267
rect 3433 4233 3467 4267
rect 3467 4233 3476 4267
rect 3424 4224 3476 4233
rect 3884 4224 3936 4276
rect 4436 4224 4488 4276
rect 2964 4088 3016 4140
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 3976 4088 4028 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 5448 4224 5500 4276
rect 5540 4224 5592 4276
rect 6736 4224 6788 4276
rect 8484 4224 8536 4276
rect 5264 4156 5316 4208
rect 4896 4088 4948 4140
rect 9588 4267 9640 4276
rect 9588 4233 9597 4267
rect 9597 4233 9631 4267
rect 9631 4233 9640 4267
rect 9588 4224 9640 4233
rect 9496 4156 9548 4208
rect 10048 4224 10100 4276
rect 11336 4224 11388 4276
rect 6920 4088 6972 4140
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8300 4088 8352 4140
rect 3976 3884 4028 3936
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 4344 3884 4396 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 9956 4131 10008 4140
rect 9956 4097 9990 4131
rect 9990 4097 10008 4131
rect 9956 4088 10008 4097
rect 11612 4088 11664 4140
rect 12164 4088 12216 4140
rect 9220 4020 9272 4072
rect 7104 3884 7156 3936
rect 7656 3884 7708 3936
rect 8668 3952 8720 4004
rect 8484 3884 8536 3936
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9128 3884 9180 3936
rect 11704 3884 11756 3936
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 3792 3680 3844 3732
rect 4068 3680 4120 3732
rect 4896 3680 4948 3732
rect 5816 3680 5868 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 13176 3680 13228 3732
rect 3516 3612 3568 3664
rect 2320 3476 2372 3528
rect 3700 3408 3752 3460
rect 4252 3612 4304 3664
rect 4620 3544 4672 3596
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 2320 3340 2372 3392
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 4712 3340 4764 3392
rect 5356 3612 5408 3664
rect 5264 3544 5316 3596
rect 5448 3476 5500 3528
rect 5632 3476 5684 3528
rect 6276 3476 6328 3528
rect 8484 3544 8536 3596
rect 9956 3544 10008 3596
rect 7104 3476 7156 3528
rect 7656 3519 7708 3528
rect 7656 3485 7690 3519
rect 7690 3485 7708 3519
rect 7656 3476 7708 3485
rect 12164 3476 12216 3528
rect 6552 3408 6604 3460
rect 13452 3408 13504 3460
rect 5632 3383 5684 3392
rect 5632 3349 5641 3383
rect 5641 3349 5675 3383
rect 5675 3349 5684 3383
rect 5632 3340 5684 3349
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 4918 3238 4970 3290
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 5238 3238 5290 3290
rect 10918 3238 10970 3290
rect 10982 3238 11034 3290
rect 11046 3238 11098 3290
rect 11110 3238 11162 3290
rect 11174 3238 11226 3290
rect 11238 3238 11290 3290
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5448 3136 5500 3188
rect 6000 3136 6052 3188
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2320 3000 2372 3052
rect 3792 3000 3844 3052
rect 6276 3000 6328 3052
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 7104 3136 7156 3188
rect 7380 3136 7432 3188
rect 9036 3136 9088 3188
rect 8576 3000 8628 3052
rect 12164 3000 12216 3052
rect 8392 2864 8444 2916
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 2964 2796 3016 2848
rect 5540 2796 5592 2848
rect 9220 2796 9272 2848
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 8484 2592 8536 2644
rect 9496 2592 9548 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 8760 2524 8812 2576
rect 9312 2524 9364 2576
rect 2872 2456 2924 2508
rect 5632 2456 5684 2508
rect 1676 2388 1728 2440
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 5540 2388 5592 2440
rect 5448 2320 5500 2372
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10600 2388 10652 2440
rect 11704 2388 11756 2440
rect 13360 2388 13412 2440
rect 14096 2388 14148 2440
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 9220 2320 9272 2372
rect 940 2252 992 2304
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 4620 2295 4672 2304
rect 4620 2261 4629 2295
rect 4629 2261 4663 2295
rect 4663 2261 4672 2295
rect 4620 2252 4672 2261
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 11796 2295 11848 2304
rect 11796 2261 11805 2295
rect 11805 2261 11839 2295
rect 11839 2261 11848 2295
rect 11796 2252 11848 2261
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 4918 2150 4970 2202
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 5238 2150 5290 2202
rect 10918 2150 10970 2202
rect 10982 2150 11034 2202
rect 11046 2150 11098 2202
rect 11110 2150 11162 2202
rect 11174 2150 11226 2202
rect 11238 2150 11290 2202
<< metal2 >>
rect 938 16435 994 17235
rect 1950 16538 2006 17235
rect 2962 16538 3018 17235
rect 1950 16510 2360 16538
rect 1950 16435 2006 16510
rect 952 14618 980 16435
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2332 14618 2360 16510
rect 2962 16510 3096 16538
rect 2962 16435 3018 16510
rect 3068 14618 3096 16510
rect 3974 16435 4030 17235
rect 4986 16538 5042 17235
rect 4986 16510 5120 16538
rect 4986 16435 5042 16510
rect 3988 14618 4016 16435
rect 5092 14618 5120 16510
rect 5998 16435 6054 17235
rect 7010 16435 7066 17235
rect 8022 16538 8078 17235
rect 7852 16510 8078 16538
rect 6012 14618 6040 16435
rect 7024 14618 7052 16435
rect 7852 14618 7880 16510
rect 8022 16435 8078 16510
rect 9034 16435 9090 17235
rect 10046 16435 10102 17235
rect 11058 16435 11114 17235
rect 12070 16435 12126 17235
rect 13082 16435 13138 17235
rect 14094 16435 14150 17235
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 9048 14618 9076 16435
rect 940 14612 992 14618
rect 940 14554 992 14560
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 1596 9178 1624 14350
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2148 12986 2176 13194
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11218 1716 12038
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1780 11354 1808 11698
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 2332 11354 2360 12786
rect 2700 12782 2728 13262
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11898 2544 12106
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2608 11354 2636 12038
rect 2700 11830 2728 12718
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 2700 10996 2728 11766
rect 2792 11558 2820 14350
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2884 13190 2912 13874
rect 2976 13190 3004 13874
rect 3252 13818 3280 14350
rect 3528 13938 3556 14486
rect 4252 14408 4304 14414
rect 4172 14368 4252 14396
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3160 13790 3280 13818
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2884 12986 2912 13126
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2884 11694 2912 12922
rect 2976 12306 3004 13126
rect 3068 12322 3096 13398
rect 3160 12434 3188 13790
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 12866 3280 13670
rect 3422 13424 3478 13433
rect 3344 13382 3422 13410
rect 3344 13326 3372 13382
rect 3422 13359 3478 13368
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3252 12850 3372 12866
rect 3252 12844 3384 12850
rect 3252 12838 3332 12844
rect 3332 12786 3384 12792
rect 3160 12406 3372 12434
rect 3344 12322 3372 12406
rect 2964 12300 3016 12306
rect 3068 12294 3188 12322
rect 3344 12294 3464 12322
rect 2964 12242 3016 12248
rect 3160 12238 3188 12294
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2884 11014 2912 11630
rect 3068 11218 3096 12038
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2872 11008 2924 11014
rect 2700 10968 2820 10996
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 2792 9654 2820 10968
rect 2872 10950 2924 10956
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1596 8498 1624 9114
rect 2792 8974 2820 9590
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1688 7954 1716 8910
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 2792 8498 2820 8910
rect 2884 8838 2912 10950
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2976 9178 3004 9454
rect 3068 9178 3096 9454
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2136 8424 2188 8430
rect 2134 8392 2136 8401
rect 2872 8424 2924 8430
rect 2188 8392 2190 8401
rect 2872 8366 2924 8372
rect 2134 8327 2190 8336
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2884 6866 2912 8366
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 7750 3004 8298
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6322 3004 6666
rect 3068 6458 3096 6734
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 2446 1716 6054
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 2976 5914 3004 6258
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 5234 1808 5510
rect 2332 5234 2360 5646
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2976 5370 3004 5578
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 2332 3534 2360 5170
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2320 3528 2372 3534
rect 2240 3488 2320 3516
rect 2240 3058 2268 3488
rect 2320 3470 2372 3476
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3058 2360 3334
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 2884 2514 2912 4966
rect 3160 4146 3188 12174
rect 3252 11830 3280 12174
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3252 11082 3280 11766
rect 3344 11694 3372 12038
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3344 11286 3372 11630
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 9450 3280 11018
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 8974 3280 9114
rect 3344 9110 3372 11222
rect 3436 10690 3464 12294
rect 3528 12102 3556 13874
rect 3712 13462 3740 14282
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3712 11898 3740 12310
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 10810 3648 11630
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3436 10662 3648 10690
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3344 8974 3372 9046
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3252 8838 3280 8910
rect 3436 8838 3464 9522
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 7954 3464 8774
rect 3528 8022 3556 9454
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3620 7750 3648 10662
rect 3804 9058 3832 13874
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13530 4016 13670
rect 4080 13530 4108 13874
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12986 3924 13126
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12640 4028 12646
rect 4028 12600 4108 12628
rect 3976 12582 4028 12588
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3988 10062 4016 11222
rect 4080 11132 4108 12600
rect 4172 11200 4200 14368
rect 4252 14350 4304 14356
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 4916 14172 5292 14181
rect 4972 14170 4996 14172
rect 5052 14170 5076 14172
rect 5132 14170 5156 14172
rect 5212 14170 5236 14172
rect 4972 14118 4982 14170
rect 5226 14118 5236 14170
rect 4972 14116 4996 14118
rect 5052 14116 5076 14118
rect 5132 14116 5156 14118
rect 5212 14116 5236 14118
rect 4916 14107 5292 14116
rect 5368 14006 5396 14350
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 4448 13433 4476 13942
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4434 13424 4490 13433
rect 4434 13359 4490 13368
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11778 4292 12106
rect 4448 11898 4476 13359
rect 4540 12986 4568 13874
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4816 12986 4844 13738
rect 5460 13546 5488 14486
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 5368 13518 5488 13546
rect 5644 13530 5672 14214
rect 6932 14074 6960 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7760 14006 7788 14350
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 7104 14000 7156 14006
rect 6748 13948 7104 13954
rect 6748 13942 7156 13948
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 6748 13938 7144 13942
rect 6736 13932 7144 13938
rect 6788 13926 7144 13932
rect 7196 13932 7248 13938
rect 6736 13874 6788 13880
rect 7196 13874 7248 13880
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 5632 13524 5684 13530
rect 5368 13258 5396 13518
rect 5632 13466 5684 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 6182 13424 6238 13433
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 4916 13084 5292 13093
rect 4972 13082 4996 13084
rect 5052 13082 5076 13084
rect 5132 13082 5156 13084
rect 5212 13082 5236 13084
rect 4972 13030 4982 13082
rect 5226 13030 5236 13082
rect 4972 13028 4996 13030
rect 5052 13028 5076 13030
rect 5132 13028 5156 13030
rect 5212 13028 5236 13030
rect 4916 13019 5292 13028
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4540 12866 4568 12922
rect 5264 12912 5316 12918
rect 4540 12838 4936 12866
rect 5264 12854 5316 12860
rect 4908 12434 4936 12838
rect 5276 12714 5304 12854
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 4540 12406 4936 12434
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4434 11792 4490 11801
rect 4264 11750 4384 11778
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4264 11558 4292 11630
rect 4252 11552 4304 11558
rect 4250 11520 4252 11529
rect 4304 11520 4306 11529
rect 4250 11455 4306 11464
rect 4356 11354 4384 11750
rect 4434 11727 4436 11736
rect 4488 11727 4490 11736
rect 4436 11698 4488 11704
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4172 11172 4292 11200
rect 4080 11104 4200 11132
rect 4172 11014 4200 11104
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4080 10810 4108 10950
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4172 10674 4200 10950
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4264 9674 4292 11172
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10742 4384 11086
rect 4540 10996 4568 12406
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4448 10968 4568 10996
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4172 9646 4292 9674
rect 4356 9654 4384 9862
rect 4344 9648 4396 9654
rect 4172 9586 4200 9646
rect 4344 9590 4396 9596
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3712 9030 3832 9058
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6458 3280 6598
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3344 5370 3372 5850
rect 3620 5778 3648 6122
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3712 5642 3740 9030
rect 3896 8974 3924 9454
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 8974 4016 9318
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3896 8838 3924 8910
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3804 7818 3832 8774
rect 4264 8634 4292 9114
rect 3976 8628 4028 8634
rect 4252 8628 4304 8634
rect 4028 8588 4200 8616
rect 3976 8570 4028 8576
rect 4172 8022 4200 8588
rect 4252 8570 4304 8576
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 8090 4292 8230
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4080 7834 4108 7958
rect 3792 7812 3844 7818
rect 4080 7806 4200 7834
rect 3792 7754 3844 7760
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3608 5568 3660 5574
rect 3804 5556 3832 6394
rect 3988 6322 4016 6802
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5914 3924 6054
rect 4080 5914 4108 6258
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3884 5568 3936 5574
rect 3804 5528 3884 5556
rect 3608 5510 3660 5516
rect 3884 5510 3936 5516
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3436 4282 3464 4558
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 2976 2854 3004 4082
rect 3528 3670 3556 4082
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 3620 2446 3648 5510
rect 3896 5370 3924 5510
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3896 4486 3924 5306
rect 3988 5234 4016 5714
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3804 3738 3832 4422
rect 3896 4282 3924 4422
rect 3988 4321 4016 5170
rect 4172 4554 4200 7806
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3974 4312 4030 4321
rect 3884 4276 3936 4282
rect 3974 4247 4030 4256
rect 3884 4218 3936 4224
rect 3988 4146 4016 4247
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3942 4016 4082
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3738 4108 3878
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4264 3670 4292 7754
rect 4448 6916 4476 10968
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4540 8906 4568 10746
rect 4632 10674 4660 12038
rect 4724 11694 4752 12310
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4816 11812 4844 12242
rect 5368 12102 5396 12582
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 4916 11996 5292 12005
rect 4972 11994 4996 11996
rect 5052 11994 5076 11996
rect 5132 11994 5156 11996
rect 5212 11994 5236 11996
rect 4972 11942 4982 11994
rect 5226 11942 5236 11994
rect 4972 11940 4996 11942
rect 5052 11940 5076 11942
rect 5132 11940 5156 11942
rect 5212 11940 5236 11942
rect 4916 11931 5292 11940
rect 5368 11898 5396 12038
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 4896 11824 4948 11830
rect 4816 11784 4896 11812
rect 4896 11766 4948 11772
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11540 4844 11630
rect 4724 11512 4844 11540
rect 4724 11150 4752 11512
rect 5000 11393 5028 11766
rect 5080 11688 5132 11694
rect 5078 11656 5080 11665
rect 5132 11656 5134 11665
rect 5078 11591 5134 11600
rect 4986 11384 5042 11393
rect 5184 11354 5212 11834
rect 5354 11384 5410 11393
rect 4986 11319 5042 11328
rect 5172 11348 5224 11354
rect 5354 11319 5410 11328
rect 5172 11290 5224 11296
rect 4896 11280 4948 11286
rect 4948 11240 5120 11268
rect 4896 11222 4948 11228
rect 5092 11150 5120 11240
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4896 11144 4948 11150
rect 5080 11144 5132 11150
rect 4986 11112 5042 11121
rect 4948 11092 4986 11098
rect 4896 11086 4986 11092
rect 4908 11070 4986 11086
rect 5080 11086 5132 11092
rect 4986 11047 5042 11056
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 9178 4660 10406
rect 4724 10266 4752 10950
rect 4816 10538 4844 10950
rect 4916 10908 5292 10917
rect 4972 10906 4996 10908
rect 5052 10906 5076 10908
rect 5132 10906 5156 10908
rect 5212 10906 5236 10908
rect 4972 10854 4982 10906
rect 5226 10854 5236 10906
rect 4972 10852 4996 10854
rect 5052 10852 5076 10854
rect 5132 10852 5156 10854
rect 5212 10852 5236 10854
rect 4916 10843 5292 10852
rect 5368 10810 5396 11319
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4816 9722 4844 10474
rect 4908 10198 4936 10610
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4916 9820 5292 9829
rect 4972 9818 4996 9820
rect 5052 9818 5076 9820
rect 5132 9818 5156 9820
rect 5212 9818 5236 9820
rect 4972 9766 4982 9818
rect 5226 9766 5236 9818
rect 4972 9764 4996 9766
rect 5052 9764 5076 9766
rect 5132 9764 5156 9766
rect 5212 9764 5236 9766
rect 4916 9755 5292 9764
rect 4804 9716 4856 9722
rect 5460 9674 5488 13398
rect 6182 13359 6184 13368
rect 6236 13359 6238 13368
rect 6184 13330 6236 13336
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5736 12442 5764 13262
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5828 12442 5856 12922
rect 6288 12782 6316 13466
rect 6380 13258 6408 13466
rect 6656 13410 6684 13806
rect 6748 13530 6776 13874
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13530 6868 13806
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7208 13433 7236 13874
rect 7194 13424 7250 13433
rect 6656 13394 6776 13410
rect 6656 13388 6788 13394
rect 6656 13382 6736 13388
rect 7194 13359 7250 13368
rect 6736 13330 6788 13336
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 4804 9658 4856 9664
rect 5368 9646 5488 9674
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4540 8566 4568 8842
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 7954 4660 8434
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4724 7886 4752 9046
rect 4916 8732 5292 8741
rect 4972 8730 4996 8732
rect 5052 8730 5076 8732
rect 5132 8730 5156 8732
rect 5212 8730 5236 8732
rect 4972 8678 4982 8730
rect 5226 8678 5236 8730
rect 4972 8676 4996 8678
rect 5052 8676 5076 8678
rect 5132 8676 5156 8678
rect 5212 8676 5236 8678
rect 4916 8667 5292 8676
rect 5368 8616 5396 9646
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9042 5488 9454
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5552 8974 5580 12174
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11286 5672 11698
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 8974 5672 11086
rect 5736 10674 5764 12038
rect 5828 11558 5856 12174
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5920 11218 5948 12174
rect 6012 11830 6040 12378
rect 6000 11824 6052 11830
rect 5998 11792 6000 11801
rect 6052 11792 6054 11801
rect 5998 11727 6054 11736
rect 6012 11540 6040 11727
rect 6104 11694 6132 12378
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6012 11512 6132 11540
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 11098 6040 11154
rect 5920 11070 6040 11098
rect 5920 11014 5948 11070
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6000 11008 6052 11014
rect 6104 10985 6132 11512
rect 6196 11218 6224 12106
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6288 11234 6316 11562
rect 6380 11354 6408 13194
rect 6460 13184 6512 13190
rect 6644 13184 6696 13190
rect 6512 13144 6644 13172
rect 6460 13126 6512 13132
rect 6644 13126 6696 13132
rect 6748 12442 6776 13330
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12986 7236 13262
rect 7760 12986 7788 13942
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 8588 13190 8616 14214
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 8680 13530 8708 13874
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 9692 13326 9720 13806
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 6736 12436 6788 12442
rect 7760 12434 7788 12922
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 6736 12378 6788 12384
rect 7208 12406 7788 12434
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6184 11212 6236 11218
rect 6288 11206 6408 11234
rect 6184 11154 6236 11160
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6000 10950 6052 10956
rect 6090 10976 6146 10985
rect 6012 10674 6040 10950
rect 6090 10911 6146 10920
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10266 5856 10406
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5184 8588 5396 8616
rect 5184 8362 5212 8588
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8090 5120 8230
rect 5368 8090 5396 8298
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4356 6888 4476 6916
rect 4356 3942 4384 6888
rect 4540 6322 4568 7822
rect 4816 6798 4844 7958
rect 5460 7886 5488 7958
rect 4988 7880 5040 7886
rect 4986 7848 4988 7857
rect 5356 7880 5408 7886
rect 5040 7848 5042 7857
rect 5356 7822 5408 7828
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 4986 7783 5042 7792
rect 4916 7644 5292 7653
rect 4972 7642 4996 7644
rect 5052 7642 5076 7644
rect 5132 7642 5156 7644
rect 5212 7642 5236 7644
rect 4972 7590 4982 7642
rect 5226 7590 5236 7642
rect 4972 7588 4996 7590
rect 5052 7588 5076 7590
rect 5132 7588 5156 7590
rect 5212 7588 5236 7590
rect 4916 7579 5292 7588
rect 5368 7478 5396 7822
rect 5552 7546 5580 8910
rect 5644 8430 5672 8910
rect 5828 8634 5856 9046
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7886 5764 8230
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5644 7410 5672 7822
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4448 5370 4476 5782
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4540 5302 4568 6122
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4632 5114 4660 6054
rect 4724 5234 4752 6190
rect 4816 5574 4844 6598
rect 4916 6556 5292 6565
rect 4972 6554 4996 6556
rect 5052 6554 5076 6556
rect 5132 6554 5156 6556
rect 5212 6554 5236 6556
rect 4972 6502 4982 6554
rect 5226 6502 5236 6554
rect 4972 6500 4996 6502
rect 5052 6500 5076 6502
rect 5132 6500 5156 6502
rect 5212 6500 5236 6502
rect 4916 6491 5292 6500
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 4916 5468 5292 5477
rect 4972 5466 4996 5468
rect 5052 5466 5076 5468
rect 5132 5466 5156 5468
rect 5212 5466 5236 5468
rect 4972 5414 4982 5466
rect 5226 5414 5236 5466
rect 4972 5412 4996 5414
rect 5052 5412 5076 5414
rect 5132 5412 5156 5414
rect 5212 5412 5236 5414
rect 4916 5403 5292 5412
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5356 5160 5408 5166
rect 4632 5098 4752 5114
rect 5356 5102 5408 5108
rect 4632 5092 4764 5098
rect 4632 5086 4712 5092
rect 4712 5034 4764 5040
rect 4724 4622 4752 5034
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4434 4312 4490 4321
rect 4724 4298 4752 4558
rect 4434 4247 4436 4256
rect 4488 4247 4490 4256
rect 4540 4270 4752 4298
rect 4436 4218 4488 4224
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 4049 4476 4082
rect 4434 4040 4490 4049
rect 4434 3975 4490 3984
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4540 3618 4568 4270
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4540 3602 4660 3618
rect 4540 3596 4672 3602
rect 4540 3590 4620 3596
rect 4620 3538 4672 3544
rect 4724 3534 4752 3878
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3712 3194 3740 3402
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3804 3058 3832 3334
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4724 2774 4752 3334
rect 4816 3194 4844 4558
rect 5368 4486 5396 5102
rect 5552 4622 5580 5170
rect 5540 4616 5592 4622
rect 5460 4576 5540 4604
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 4916 4380 5292 4389
rect 4972 4378 4996 4380
rect 5052 4378 5076 4380
rect 5132 4378 5156 4380
rect 5212 4378 5236 4380
rect 4972 4326 4982 4378
rect 5226 4326 5236 4378
rect 4972 4324 4996 4326
rect 5052 4324 5076 4326
rect 5132 4324 5156 4326
rect 5212 4324 5236 4326
rect 4916 4315 5292 4324
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3738 4936 4082
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5276 3602 5304 4150
rect 5368 3670 5396 4422
rect 5460 4282 5488 4576
rect 5540 4558 5592 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4282 5580 4422
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5460 3534 5488 4218
rect 5644 3534 5672 5510
rect 5736 5234 5764 7210
rect 5828 7206 5856 8570
rect 5920 8430 5948 9590
rect 6288 9382 6316 11018
rect 6380 10810 6408 11206
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6380 9926 6408 10474
rect 6472 10062 6500 11494
rect 6564 11354 6592 11630
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6840 11234 6868 11630
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11354 6960 11562
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6918 11248 6974 11257
rect 6564 11206 6918 11234
rect 6564 11150 6592 11206
rect 6918 11183 6974 11192
rect 6552 11144 6604 11150
rect 6736 11144 6788 11150
rect 6552 11086 6604 11092
rect 6656 11092 6736 11098
rect 6788 11104 6868 11132
rect 6656 11086 6788 11092
rect 6656 11070 6776 11086
rect 6656 10742 6684 11070
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 10198 6592 10610
rect 6656 10606 6684 10678
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6748 10198 6776 10950
rect 6840 10849 6868 11104
rect 6826 10840 6882 10849
rect 6826 10775 6882 10784
rect 6826 10704 6882 10713
rect 6826 10639 6828 10648
rect 6880 10639 6882 10648
rect 6828 10610 6880 10616
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10266 6868 10406
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6380 9194 6408 9862
rect 6288 9166 6408 9194
rect 6288 8974 6316 9166
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6368 8968 6420 8974
rect 6472 8922 6500 9998
rect 6564 9586 6592 10134
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6656 9674 6684 10066
rect 6840 10062 6868 10202
rect 6932 10062 6960 11183
rect 7024 10266 7052 11494
rect 7116 11354 7144 12106
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7208 11234 7236 12406
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7654 11656 7710 11665
rect 7116 11206 7236 11234
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6656 9654 6776 9674
rect 6656 9648 6788 9654
rect 6656 9646 6736 9648
rect 6736 9590 6788 9596
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6840 9382 6868 9998
rect 6932 9518 6960 9998
rect 7116 9602 7144 11206
rect 7300 11082 7328 11630
rect 7484 11286 7512 11630
rect 7654 11591 7710 11600
rect 7840 11620 7892 11626
rect 7668 11286 7696 11591
rect 7840 11562 7892 11568
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7194 10976 7250 10985
rect 7194 10911 7250 10920
rect 7208 10266 7236 10911
rect 7300 10606 7328 11018
rect 7392 10810 7420 11018
rect 7484 10810 7512 11222
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7378 10704 7434 10713
rect 7378 10639 7434 10648
rect 7656 10668 7708 10674
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7024 9574 7144 9602
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6420 8916 6500 8922
rect 6368 8910 6500 8916
rect 6380 8894 6500 8910
rect 6932 8906 6960 9454
rect 6552 8900 6604 8906
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6196 7954 6224 8570
rect 6288 8566 6316 8774
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6380 7954 6408 8894
rect 6552 8842 6604 8848
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6000 7880 6052 7886
rect 6380 7834 6408 7890
rect 6052 7828 6408 7834
rect 6000 7822 6408 7828
rect 6012 7806 6408 7822
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6012 7410 6040 7686
rect 6104 7546 6132 7686
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5920 7002 5948 7346
rect 6472 7342 6500 8570
rect 6564 8498 6592 8842
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8634 6684 8774
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6656 7954 6684 8570
rect 6932 8498 6960 8842
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6840 7834 6868 8230
rect 6840 7806 6960 7834
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6748 7342 6776 7482
rect 6932 7410 6960 7806
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6458 6316 6734
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6472 5234 6500 7142
rect 6920 6792 6972 6798
rect 6918 6760 6920 6769
rect 6972 6760 6974 6769
rect 6918 6695 6974 6704
rect 6920 6384 6972 6390
rect 7024 6372 7052 9574
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 8294 7144 9386
rect 7208 9178 7236 10066
rect 7300 9926 7328 10542
rect 7392 10062 7420 10639
rect 7656 10610 7708 10616
rect 7668 10130 7696 10610
rect 7760 10470 7788 11290
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7852 10266 7880 11562
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 7930 11248 7986 11257
rect 7930 11183 7986 11192
rect 7944 11150 7972 11183
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8300 11144 8352 11150
rect 8588 11132 8616 13126
rect 8956 12918 8984 13126
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 9232 12782 9260 13126
rect 9784 12986 9812 13874
rect 10060 13705 10088 16435
rect 11072 14414 11100 16435
rect 12084 14414 12112 16435
rect 13096 14414 13124 16435
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 10916 14172 11292 14181
rect 10972 14170 10996 14172
rect 11052 14170 11076 14172
rect 11132 14170 11156 14172
rect 11212 14170 11236 14172
rect 10972 14118 10982 14170
rect 11226 14118 11236 14170
rect 10972 14116 10996 14118
rect 11052 14116 11076 14118
rect 11132 14116 11156 14118
rect 11212 14116 11236 14118
rect 10916 14107 11292 14116
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10152 13841 10180 13874
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 10692 13728 10744 13734
rect 10046 13696 10102 13705
rect 10692 13670 10744 13676
rect 10046 13631 10102 13640
rect 10704 13258 10732 13670
rect 10888 13274 10916 13874
rect 11348 13308 11376 14214
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11348 13280 11468 13308
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10796 13246 10916 13274
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 8680 12374 8708 12718
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8680 11762 8708 12310
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11286 8708 11494
rect 8956 11354 8984 12582
rect 9232 12238 9260 12582
rect 9508 12434 9536 12786
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9324 12406 9536 12434
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11558 9260 12174
rect 9324 12102 9352 12406
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9324 11694 9352 12038
rect 9416 11830 9444 12038
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 9232 11150 9260 11494
rect 9220 11144 9272 11150
rect 8300 11086 8352 11092
rect 8482 11112 8538 11121
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10849 7972 10950
rect 7930 10840 7986 10849
rect 7930 10775 7986 10784
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8036 10713 8064 10746
rect 8022 10704 8078 10713
rect 8312 10674 8340 11086
rect 8392 11076 8444 11082
rect 8588 11104 8708 11132
rect 8482 11047 8538 11056
rect 8392 11018 8444 11024
rect 8022 10639 8078 10648
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 7840 10260 7892 10266
rect 7760 10220 7840 10248
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7116 7886 7144 8230
rect 7208 8090 7236 9114
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7116 7478 7144 7822
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7116 6798 7144 7414
rect 7208 7002 7236 7686
rect 7300 7410 7328 9862
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8090 7420 9318
rect 7484 9178 7512 9998
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7760 8838 7788 10220
rect 7840 10202 7892 10208
rect 8404 9994 8432 11018
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 7852 9722 7880 9930
rect 8496 9926 8524 11047
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10674 8616 10950
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10062 8616 10610
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 7840 9716 7892 9722
rect 8680 9674 8708 11104
rect 9220 11086 9272 11092
rect 9034 10840 9090 10849
rect 9034 10775 9090 10784
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 7840 9658 7892 9664
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7852 8634 7880 9658
rect 8496 9646 8708 9674
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7392 7410 7420 7890
rect 7576 7546 7604 8570
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 8022 7788 8434
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7760 7410 7788 7958
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7300 6934 7328 7346
rect 7484 7290 7512 7346
rect 7392 7262 7512 7290
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6972 6344 7052 6372
rect 6920 6326 6972 6332
rect 7392 6322 7420 7262
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 6322 7512 6802
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6564 5098 6592 5578
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 5736 4622 5764 5034
rect 6656 4826 6684 5170
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 3738 5856 4558
rect 6748 4554 6776 4762
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 4916 3292 5292 3301
rect 4972 3290 4996 3292
rect 5052 3290 5076 3292
rect 5132 3290 5156 3292
rect 5212 3290 5236 3292
rect 4972 3238 4982 3290
rect 5226 3238 5236 3290
rect 4972 3236 4996 3238
rect 5052 3236 5076 3238
rect 5132 3236 5156 3238
rect 5212 3236 5236 3238
rect 4916 3227 5292 3236
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 4724 2746 4844 2774
rect 4816 2446 4844 2746
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5460 2378 5488 3130
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2446 5580 2790
rect 5644 2514 5672 3334
rect 6012 3194 6040 4422
rect 6748 4282 6776 4490
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6932 4146 6960 5238
rect 7116 5234 7144 6054
rect 7392 5914 7420 6258
rect 7668 6186 7696 7278
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7760 5846 7788 6938
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5710 7880 8570
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8404 7750 8432 8026
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7478 8432 7686
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 7290 8340 7346
rect 8312 7262 8432 7290
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8036 6322 8064 6666
rect 8312 6322 8340 6734
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8312 6118 8340 6258
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8404 5914 8432 7262
rect 8496 6254 8524 9646
rect 8772 8974 8800 10406
rect 8956 10266 8984 10610
rect 9048 10266 9076 10775
rect 9416 10674 9444 11766
rect 9600 11762 9628 12038
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9600 10538 9628 11698
rect 9692 11558 9720 12174
rect 9784 12152 9812 12582
rect 9876 12442 9904 12922
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9968 12238 9996 12378
rect 10322 12336 10378 12345
rect 10322 12271 10378 12280
rect 9956 12232 10008 12238
rect 10230 12200 10286 12209
rect 9956 12174 10008 12180
rect 9864 12164 9916 12170
rect 9784 12124 9864 12152
rect 9864 12106 9916 12112
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10152 12158 10230 12186
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9784 11370 9812 11766
rect 9692 11342 9812 11370
rect 9692 10538 9720 11342
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9404 10464 9456 10470
rect 9692 10441 9720 10474
rect 9404 10406 9456 10412
rect 9678 10432 9734 10441
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9048 9586 9076 9862
rect 9140 9722 9168 9862
rect 9416 9722 9444 10406
rect 9678 10367 9734 10376
rect 9692 9738 9720 10367
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9508 9710 9720 9738
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8634 8800 8910
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7857 8708 7890
rect 8956 7886 8984 9318
rect 9140 8974 9168 9386
rect 9416 9178 9444 9658
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9310 8392 9366 8401
rect 9508 8378 9536 9710
rect 9678 9616 9734 9625
rect 9588 9580 9640 9586
rect 9784 9586 9812 10746
rect 9678 9551 9680 9560
rect 9588 9522 9640 9528
rect 9732 9551 9734 9560
rect 9772 9580 9824 9586
rect 9680 9522 9732 9528
rect 9772 9522 9824 9528
rect 9600 9178 9628 9522
rect 9876 9489 9904 12106
rect 10060 11762 10088 12106
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11257 9996 11494
rect 9954 11248 10010 11257
rect 9954 11183 10010 11192
rect 9862 9480 9918 9489
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9772 9444 9824 9450
rect 9862 9415 9918 9424
rect 9772 9386 9824 9392
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 8838 9720 9386
rect 9784 9217 9812 9386
rect 9770 9208 9826 9217
rect 9770 9143 9826 9152
rect 9770 9072 9826 9081
rect 9770 9007 9772 9016
rect 9824 9007 9826 9016
rect 9772 8978 9824 8984
rect 9876 8974 9904 9415
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9784 8430 9812 8842
rect 9876 8498 9904 8910
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9366 8350 9536 8378
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9310 8327 9366 8336
rect 8944 7880 8996 7886
rect 8666 7848 8722 7857
rect 8944 7822 8996 7828
rect 8666 7783 8722 7792
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8588 6390 8616 7210
rect 8680 6934 8708 7482
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6662 8800 6734
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8772 6322 8800 6598
rect 8956 6458 8984 7822
rect 9324 7546 9352 8327
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8022 9812 8230
rect 9968 8072 9996 11183
rect 10060 10742 10088 11698
rect 10152 10826 10180 12158
rect 10230 12135 10286 12144
rect 10336 11898 10364 12271
rect 10428 12238 10456 12718
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10336 11082 10364 11698
rect 10428 11558 10456 12174
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10152 10798 10456 10826
rect 10048 10736 10100 10742
rect 10100 10696 10272 10724
rect 10048 10678 10100 10684
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10060 10169 10088 10542
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 9722 10088 9930
rect 10152 9722 10180 10406
rect 10244 9722 10272 10696
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10244 9500 10272 9658
rect 10152 9472 10272 9500
rect 10152 9466 10180 9472
rect 10060 9438 10180 9466
rect 10060 8090 10088 9438
rect 10336 8956 10364 10406
rect 10428 9586 10456 10798
rect 10520 9722 10548 12174
rect 10612 12170 10640 12854
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10612 11762 10640 12106
rect 10704 11898 10732 12174
rect 10796 11898 10824 13246
rect 10916 13084 11292 13093
rect 10972 13082 10996 13084
rect 11052 13082 11076 13084
rect 11132 13082 11156 13084
rect 11212 13082 11236 13084
rect 10972 13030 10982 13082
rect 11226 13030 11236 13082
rect 10972 13028 10996 13030
rect 11052 13028 11076 13030
rect 11132 13028 11156 13030
rect 11212 13028 11236 13030
rect 10916 13019 11292 13028
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11244 12368 11296 12374
rect 10874 12336 10930 12345
rect 10930 12306 11008 12322
rect 11244 12310 11296 12316
rect 10930 12300 11020 12306
rect 10930 12294 10968 12300
rect 10874 12271 10930 12280
rect 10968 12242 11020 12248
rect 10876 12232 10928 12238
rect 10966 12200 11022 12209
rect 10928 12180 10966 12186
rect 10876 12174 10966 12180
rect 10888 12158 10966 12174
rect 10966 12135 11022 12144
rect 11256 12102 11284 12310
rect 11348 12238 11376 12650
rect 11440 12434 11468 13280
rect 11532 12986 11560 13874
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12986 11836 13126
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11440 12406 11560 12434
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10916 11996 11292 12005
rect 10972 11994 10996 11996
rect 11052 11994 11076 11996
rect 11132 11994 11156 11996
rect 11212 11994 11236 11996
rect 10972 11942 10982 11994
rect 11226 11942 11236 11994
rect 10972 11940 10996 11942
rect 11052 11940 11076 11942
rect 11132 11940 11156 11942
rect 11212 11940 11236 11942
rect 10916 11931 11292 11940
rect 11348 11898 11376 12174
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11354 10640 11698
rect 10888 11676 10916 11834
rect 10968 11756 11020 11762
rect 11244 11756 11296 11762
rect 10968 11698 11020 11704
rect 11164 11716 11244 11744
rect 10704 11648 10916 11676
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10441 10640 10610
rect 10704 10577 10732 11648
rect 10980 11558 11008 11698
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11370 11100 11494
rect 11164 11393 11192 11716
rect 11244 11698 11296 11704
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11256 11529 11284 11562
rect 11242 11520 11298 11529
rect 11242 11455 11298 11464
rect 10980 11342 11100 11370
rect 11150 11384 11206 11393
rect 10980 11150 11008 11342
rect 11150 11319 11206 11328
rect 11256 11286 11284 11455
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11348 11218 11376 11562
rect 11440 11354 11468 12174
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11426 11248 11482 11257
rect 11336 11212 11388 11218
rect 11426 11183 11482 11192
rect 11336 11154 11388 11160
rect 11440 11150 11468 11183
rect 10968 11144 11020 11150
rect 10782 11112 10838 11121
rect 10968 11086 11020 11092
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 10782 11047 10838 11056
rect 10796 10674 10824 11047
rect 10980 11014 11008 11086
rect 10968 11008 11020 11014
rect 11256 10996 11284 11086
rect 11256 10968 11468 10996
rect 10968 10950 11020 10956
rect 10916 10908 11292 10917
rect 10972 10906 10996 10908
rect 11052 10906 11076 10908
rect 11132 10906 11156 10908
rect 11212 10906 11236 10908
rect 10972 10854 10982 10906
rect 11226 10854 11236 10906
rect 10972 10852 10996 10854
rect 11052 10852 11076 10854
rect 11132 10852 11156 10854
rect 11212 10852 11236 10854
rect 10916 10843 11292 10852
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11072 10577 11100 10610
rect 10690 10568 10746 10577
rect 11058 10568 11114 10577
rect 10690 10503 10746 10512
rect 10784 10532 10836 10538
rect 11058 10503 11114 10512
rect 10784 10474 10836 10480
rect 10796 10441 10824 10474
rect 10598 10432 10654 10441
rect 10598 10367 10654 10376
rect 10782 10432 10838 10441
rect 10782 10367 10838 10376
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10416 9376 10468 9382
rect 10520 9353 10548 9658
rect 10416 9318 10468 9324
rect 10506 9344 10562 9353
rect 10428 9178 10456 9318
rect 10506 9279 10562 9288
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10416 8968 10468 8974
rect 10230 8936 10286 8945
rect 10336 8928 10416 8956
rect 10416 8910 10468 8916
rect 10230 8871 10286 8880
rect 10244 8294 10272 8871
rect 10520 8838 10548 9279
rect 10612 9042 10640 10367
rect 10690 10160 10746 10169
rect 10690 10095 10746 10104
rect 10704 10062 10732 10095
rect 11072 10062 11100 10503
rect 11164 10470 11192 10746
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11256 9926 11284 10678
rect 11334 10568 11390 10577
rect 11334 10503 11390 10512
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 10704 9636 10732 9862
rect 10916 9820 11292 9829
rect 10972 9818 10996 9820
rect 11052 9818 11076 9820
rect 11132 9818 11156 9820
rect 11212 9818 11236 9820
rect 10972 9766 10982 9818
rect 11226 9766 11236 9818
rect 10972 9764 10996 9766
rect 11052 9764 11076 9766
rect 11132 9764 11156 9766
rect 11212 9764 11236 9766
rect 10916 9755 11292 9764
rect 11244 9648 11296 9654
rect 10704 9608 11192 9636
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10704 9217 10732 9454
rect 10690 9208 10746 9217
rect 10888 9178 10916 9454
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10690 9143 10746 9152
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10600 9036 10652 9042
rect 10876 9036 10928 9042
rect 10600 8978 10652 8984
rect 10796 8996 10876 9024
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10508 8832 10560 8838
rect 10612 8809 10640 8842
rect 10508 8774 10560 8780
rect 10598 8800 10654 8809
rect 10520 8616 10548 8774
rect 10598 8735 10654 8744
rect 10520 8588 10640 8616
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 9876 8044 9996 8072
rect 10048 8084 10100 8090
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9508 7002 9536 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9048 6390 9076 6938
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9402 6760 9458 6769
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9048 6254 9076 6326
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9140 6186 9168 6666
rect 9324 6662 9352 6734
rect 9784 6730 9812 7686
rect 9876 7002 9904 8044
rect 10048 8026 10100 8032
rect 9954 7984 10010 7993
rect 9954 7919 10010 7928
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9402 6695 9458 6704
rect 9680 6724 9732 6730
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7392 4690 7420 5306
rect 8312 5302 8340 5714
rect 8404 5302 8432 5850
rect 8496 5710 8524 6054
rect 9140 5846 9168 6122
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8496 5234 8524 5646
rect 9048 5370 9076 5646
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9140 5234 9168 5782
rect 9232 5710 9260 6326
rect 9324 6186 9352 6598
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9324 5710 9352 6122
rect 9416 6118 9444 6695
rect 9680 6666 9732 6672
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9692 6361 9720 6666
rect 9678 6352 9734 6361
rect 9588 6316 9640 6322
rect 9678 6287 9734 6296
rect 9588 6258 9640 6264
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9600 5846 9628 6258
rect 9784 6202 9812 6666
rect 9692 6174 9812 6202
rect 9588 5840 9640 5846
rect 9508 5800 9588 5828
rect 9508 5710 9536 5800
rect 9588 5782 9640 5788
rect 9692 5778 9720 6174
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5817 9812 6054
rect 9770 5808 9826 5817
rect 9680 5772 9732 5778
rect 9770 5743 9826 5752
rect 9680 5714 9732 5720
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9312 5704 9364 5710
rect 9496 5704 9548 5710
rect 9364 5664 9444 5692
rect 9312 5646 9364 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9324 5030 9352 5510
rect 9416 5370 9444 5664
rect 9496 5646 9548 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 3534 7144 3878
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6288 3058 6316 3470
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6564 3194 6592 3402
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 3194 7144 3334
rect 7392 3194 7420 4626
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8128 4146 8156 4422
rect 8312 4146 8340 4422
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3534 7696 3878
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 8404 2922 8432 4626
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 4282 8524 4490
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3602 8524 3878
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3058 8616 4558
rect 8680 4010 8708 4966
rect 9140 4690 9168 4966
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9324 4622 9352 4966
rect 9508 4826 9536 5238
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9692 4758 9720 5510
rect 9876 5234 9904 6938
rect 9968 6934 9996 7919
rect 10520 7886 10548 8434
rect 10612 8362 10640 8588
rect 10796 8498 10824 8996
rect 10876 8978 10928 8984
rect 10980 8974 11008 9318
rect 11060 9104 11112 9110
rect 11058 9072 11060 9081
rect 11112 9072 11114 9081
rect 11058 9007 11114 9016
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11164 8820 11192 9608
rect 11244 9590 11296 9596
rect 11256 9042 11284 9590
rect 11348 9042 11376 10503
rect 11440 10470 11468 10968
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 9586 11468 10406
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8945 11376 8978
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11164 8792 11376 8820
rect 10916 8732 11292 8741
rect 10972 8730 10996 8732
rect 11052 8730 11076 8732
rect 11132 8730 11156 8732
rect 11212 8730 11236 8732
rect 10972 8678 10982 8730
rect 11226 8678 11236 8730
rect 10972 8676 10996 8678
rect 11052 8676 11076 8678
rect 11132 8676 11156 8678
rect 11212 8676 11236 8678
rect 10916 8667 11292 8676
rect 11150 8528 11206 8537
rect 10784 8492 10836 8498
rect 11150 8463 11152 8472
rect 10784 8434 10836 8440
rect 11204 8463 11206 8472
rect 11152 8434 11204 8440
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10612 8090 10640 8298
rect 10796 8090 10824 8434
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10888 7886 10916 8366
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7206 10088 7686
rect 10916 7644 11292 7653
rect 10972 7642 10996 7644
rect 11052 7642 11076 7644
rect 11132 7642 11156 7644
rect 11212 7642 11236 7644
rect 10972 7590 10982 7642
rect 11226 7590 11236 7642
rect 10972 7588 10996 7590
rect 11052 7588 11076 7590
rect 11132 7588 11156 7590
rect 11212 7588 11236 7590
rect 10916 7579 11292 7588
rect 11348 7290 11376 8792
rect 11440 8634 11468 9522
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11532 7546 11560 12406
rect 11624 12306 11652 12786
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12374 11836 12718
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11624 11898 11652 12242
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11286 11652 11562
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10606 11652 10950
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11716 10266 11744 12242
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11898 11836 12038
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11808 10577 11836 11834
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11716 10130 11744 10202
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11716 9722 11744 10066
rect 11808 9722 11836 10066
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11900 9602 11928 14214
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12084 12238 12112 13262
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12162 12200 12218 12209
rect 12162 12135 12218 12144
rect 12256 12164 12308 12170
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11992 11898 12020 12038
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11808 9586 11928 9602
rect 11796 9580 11928 9586
rect 11848 9574 11928 9580
rect 11796 9522 11848 9528
rect 11610 9480 11666 9489
rect 11666 9438 11744 9466
rect 11610 9415 11666 9424
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11624 8498 11652 9143
rect 11716 9042 11744 9438
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11532 7426 11560 7482
rect 11440 7410 11560 7426
rect 11428 7404 11560 7410
rect 11480 7398 11560 7404
rect 11428 7346 11480 7352
rect 11520 7336 11572 7342
rect 11348 7262 11468 7290
rect 11520 7278 11572 7284
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9968 4842 9996 6870
rect 10244 6866 10272 7142
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 6322 10088 6394
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 10060 5710 10088 6151
rect 10152 5914 10180 6666
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10244 5234 10272 6802
rect 10784 6792 10836 6798
rect 10704 6752 10784 6780
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9876 4814 9996 4842
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 4282 9628 4490
rect 9876 4486 9904 4814
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 8496 2650 8524 2858
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8772 2582 8800 3334
rect 9048 3194 9076 3878
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 9140 2378 9168 3878
rect 9232 2854 9260 4014
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2378 9260 2790
rect 9508 2650 9536 4150
rect 9968 4146 9996 4694
rect 10060 4282 10088 4966
rect 10704 4826 10732 6752
rect 10784 6734 10836 6740
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 5370 10824 6598
rect 10916 6556 11292 6565
rect 10972 6554 10996 6556
rect 11052 6554 11076 6556
rect 11132 6554 11156 6556
rect 11212 6554 11236 6556
rect 10972 6502 10982 6554
rect 11226 6502 11236 6554
rect 10972 6500 10996 6502
rect 11052 6500 11076 6502
rect 11132 6500 11156 6502
rect 11212 6500 11236 6502
rect 10916 6491 11292 6500
rect 11348 6458 11376 6666
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 6390 11468 7262
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10980 6118 11008 6258
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5914 11008 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10916 5468 11292 5477
rect 10972 5466 10996 5468
rect 11052 5466 11076 5468
rect 11132 5466 11156 5468
rect 11212 5466 11236 5468
rect 10972 5414 10982 5466
rect 11226 5414 11236 5466
rect 10972 5412 10996 5414
rect 11052 5412 11076 5414
rect 11132 5412 11156 5414
rect 11212 5412 11236 5414
rect 10916 5403 11292 5412
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 11348 5234 11376 6258
rect 11532 5370 11560 7278
rect 11624 6798 11652 8434
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 6798 11744 7346
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11808 5370 11836 9522
rect 11992 8974 12020 11222
rect 12084 11150 12112 12038
rect 12176 11898 12204 12135
rect 12256 12106 12308 12112
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12268 11830 12296 12106
rect 12256 11824 12308 11830
rect 12162 11792 12218 11801
rect 12256 11766 12308 11772
rect 12162 11727 12164 11736
rect 12216 11727 12218 11736
rect 12164 11698 12216 11704
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10810 12112 10950
rect 12176 10810 12204 11494
rect 12360 11150 12388 12582
rect 12452 11898 12480 12650
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11529 12572 12650
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11830 12664 12038
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12728 11393 12756 12582
rect 12714 11384 12770 11393
rect 12714 11319 12770 11328
rect 12348 11144 12400 11150
rect 12346 11112 12348 11121
rect 13360 11144 13412 11150
rect 12400 11112 12402 11121
rect 13360 11086 13412 11092
rect 12346 11047 12402 11056
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12176 10554 12204 10746
rect 12072 10532 12124 10538
rect 12176 10526 12296 10554
rect 12072 10474 12124 10480
rect 12084 10441 12112 10474
rect 12164 10464 12216 10470
rect 12070 10432 12126 10441
rect 12164 10406 12216 10412
rect 12070 10367 12126 10376
rect 12176 10062 12204 10406
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12268 9926 12296 10526
rect 12544 10198 12572 10950
rect 12728 10742 12756 10950
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 9042 12112 9522
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12176 8634 12204 8842
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8498 12296 9862
rect 12544 8906 12572 10134
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12636 8634 12664 9930
rect 12728 9178 12756 10678
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 10062 13032 10610
rect 13188 10606 13216 10950
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 13004 8838 13032 9998
rect 13372 9450 13400 11086
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 13004 8498 13032 8774
rect 13372 8498 13400 9386
rect 14108 8566 14136 16435
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11900 6798 11928 7346
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12072 5840 12124 5846
rect 12070 5808 12072 5817
rect 12124 5808 12126 5817
rect 12070 5743 12126 5752
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 12176 5234 12204 5646
rect 12360 5302 12388 6598
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13372 5710 13400 6190
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4826 11100 4966
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10916 4380 11292 4389
rect 10972 4378 10996 4380
rect 11052 4378 11076 4380
rect 11132 4378 11156 4380
rect 11212 4378 11236 4380
rect 10972 4326 10982 4378
rect 11226 4326 11236 4378
rect 10972 4324 10996 4326
rect 11052 4324 11076 4326
rect 11132 4324 11156 4326
rect 11212 4324 11236 4326
rect 10916 4315 11292 4324
rect 11348 4282 11376 5170
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11624 4146 11652 4422
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 10138 4040 10194 4049
rect 10138 3975 10194 3984
rect 10152 3738 10180 3975
rect 11716 3942 11744 5170
rect 12176 4146 12204 5170
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 940 2304 992 2310
rect 2228 2304 2280 2310
rect 940 2246 992 2252
rect 2148 2264 2228 2292
rect 952 800 980 2246
rect 2148 800 2176 2264
rect 3424 2304 3476 2310
rect 2228 2246 2280 2252
rect 3344 2264 3424 2292
rect 3344 800 3372 2264
rect 4620 2304 4672 2310
rect 3424 2246 3476 2252
rect 4540 2264 4620 2292
rect 4540 800 4568 2264
rect 5816 2304 5868 2310
rect 4620 2246 4672 2252
rect 5736 2264 5816 2292
rect 4916 2204 5292 2213
rect 4972 2202 4996 2204
rect 5052 2202 5076 2204
rect 5132 2202 5156 2204
rect 5212 2202 5236 2204
rect 4972 2150 4982 2202
rect 5226 2150 5236 2202
rect 4972 2148 4996 2150
rect 5052 2148 5076 2150
rect 5132 2148 5156 2150
rect 5212 2148 5236 2150
rect 4916 2139 5292 2148
rect 5736 800 5764 2264
rect 5816 2246 5868 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 7024 1170 7052 2246
rect 8220 1170 8248 2246
rect 6932 1142 7052 1170
rect 8128 1142 8248 1170
rect 6932 800 6960 1142
rect 8128 800 8156 1142
rect 9324 800 9352 2518
rect 9968 2446 9996 3538
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 2446 10640 3334
rect 10916 3292 11292 3301
rect 10972 3290 10996 3292
rect 11052 3290 11076 3292
rect 11132 3290 11156 3292
rect 11212 3290 11236 3292
rect 10972 3238 10982 3290
rect 11226 3238 11236 3290
rect 10972 3236 10996 3238
rect 11052 3236 11076 3238
rect 11132 3236 11156 3238
rect 11212 3236 11236 3238
rect 10916 3227 11292 3236
rect 11716 2446 11744 3878
rect 12176 3534 12204 4082
rect 13188 3738 13216 5578
rect 13464 5370 13492 6734
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13464 3618 13492 5306
rect 13372 3590 13492 3618
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12176 3058 12204 3470
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 13372 2446 13400 3590
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13464 2650 13492 3402
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 10612 1170 10640 2246
rect 10916 2204 11292 2213
rect 10972 2202 10996 2204
rect 11052 2202 11076 2204
rect 11132 2202 11156 2204
rect 11212 2202 11236 2204
rect 10972 2150 10982 2202
rect 11226 2150 11236 2202
rect 10972 2148 10996 2150
rect 11052 2148 11076 2150
rect 11132 2148 11156 2150
rect 11212 2148 11236 2150
rect 10916 2139 11292 2148
rect 11808 1170 11836 2246
rect 13004 1170 13032 2246
rect 10520 1142 10640 1170
rect 11716 1142 11836 1170
rect 12912 1142 13032 1170
rect 10520 800 10548 1142
rect 11716 800 11744 1142
rect 12912 800 12940 1142
rect 14108 800 14136 2382
rect 938 0 994 800
rect 2134 0 2190 800
rect 3330 0 3386 800
rect 4526 0 4582 800
rect 5722 0 5778 800
rect 6918 0 6974 800
rect 8114 0 8170 800
rect 9310 0 9366 800
rect 10506 0 10562 800
rect 11702 0 11758 800
rect 12898 0 12954 800
rect 14094 0 14150 800
<< via2 >>
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 3422 13368 3478 13424
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 2134 8372 2136 8392
rect 2136 8372 2188 8392
rect 2188 8372 2190 8392
rect 2134 8336 2190 8372
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 4916 14170 4972 14172
rect 4996 14170 5052 14172
rect 5076 14170 5132 14172
rect 5156 14170 5212 14172
rect 5236 14170 5292 14172
rect 4916 14118 4918 14170
rect 4918 14118 4970 14170
rect 4970 14118 4972 14170
rect 4996 14118 5034 14170
rect 5034 14118 5046 14170
rect 5046 14118 5052 14170
rect 5076 14118 5098 14170
rect 5098 14118 5110 14170
rect 5110 14118 5132 14170
rect 5156 14118 5162 14170
rect 5162 14118 5174 14170
rect 5174 14118 5212 14170
rect 5236 14118 5238 14170
rect 5238 14118 5290 14170
rect 5290 14118 5292 14170
rect 4916 14116 4972 14118
rect 4996 14116 5052 14118
rect 5076 14116 5132 14118
rect 5156 14116 5212 14118
rect 5236 14116 5292 14118
rect 4434 13368 4490 13424
rect 4916 13082 4972 13084
rect 4996 13082 5052 13084
rect 5076 13082 5132 13084
rect 5156 13082 5212 13084
rect 5236 13082 5292 13084
rect 4916 13030 4918 13082
rect 4918 13030 4970 13082
rect 4970 13030 4972 13082
rect 4996 13030 5034 13082
rect 5034 13030 5046 13082
rect 5046 13030 5052 13082
rect 5076 13030 5098 13082
rect 5098 13030 5110 13082
rect 5110 13030 5132 13082
rect 5156 13030 5162 13082
rect 5162 13030 5174 13082
rect 5174 13030 5212 13082
rect 5236 13030 5238 13082
rect 5238 13030 5290 13082
rect 5290 13030 5292 13082
rect 4916 13028 4972 13030
rect 4996 13028 5052 13030
rect 5076 13028 5132 13030
rect 5156 13028 5212 13030
rect 5236 13028 5292 13030
rect 4250 11500 4252 11520
rect 4252 11500 4304 11520
rect 4304 11500 4306 11520
rect 4250 11464 4306 11500
rect 4434 11756 4490 11792
rect 4434 11736 4436 11756
rect 4436 11736 4488 11756
rect 4488 11736 4490 11756
rect 3974 4256 4030 4312
rect 4916 11994 4972 11996
rect 4996 11994 5052 11996
rect 5076 11994 5132 11996
rect 5156 11994 5212 11996
rect 5236 11994 5292 11996
rect 4916 11942 4918 11994
rect 4918 11942 4970 11994
rect 4970 11942 4972 11994
rect 4996 11942 5034 11994
rect 5034 11942 5046 11994
rect 5046 11942 5052 11994
rect 5076 11942 5098 11994
rect 5098 11942 5110 11994
rect 5110 11942 5132 11994
rect 5156 11942 5162 11994
rect 5162 11942 5174 11994
rect 5174 11942 5212 11994
rect 5236 11942 5238 11994
rect 5238 11942 5290 11994
rect 5290 11942 5292 11994
rect 4916 11940 4972 11942
rect 4996 11940 5052 11942
rect 5076 11940 5132 11942
rect 5156 11940 5212 11942
rect 5236 11940 5292 11942
rect 5078 11636 5080 11656
rect 5080 11636 5132 11656
rect 5132 11636 5134 11656
rect 5078 11600 5134 11636
rect 4986 11328 5042 11384
rect 5354 11328 5410 11384
rect 4986 11056 5042 11112
rect 4916 10906 4972 10908
rect 4996 10906 5052 10908
rect 5076 10906 5132 10908
rect 5156 10906 5212 10908
rect 5236 10906 5292 10908
rect 4916 10854 4918 10906
rect 4918 10854 4970 10906
rect 4970 10854 4972 10906
rect 4996 10854 5034 10906
rect 5034 10854 5046 10906
rect 5046 10854 5052 10906
rect 5076 10854 5098 10906
rect 5098 10854 5110 10906
rect 5110 10854 5132 10906
rect 5156 10854 5162 10906
rect 5162 10854 5174 10906
rect 5174 10854 5212 10906
rect 5236 10854 5238 10906
rect 5238 10854 5290 10906
rect 5290 10854 5292 10906
rect 4916 10852 4972 10854
rect 4996 10852 5052 10854
rect 5076 10852 5132 10854
rect 5156 10852 5212 10854
rect 5236 10852 5292 10854
rect 4916 9818 4972 9820
rect 4996 9818 5052 9820
rect 5076 9818 5132 9820
rect 5156 9818 5212 9820
rect 5236 9818 5292 9820
rect 4916 9766 4918 9818
rect 4918 9766 4970 9818
rect 4970 9766 4972 9818
rect 4996 9766 5034 9818
rect 5034 9766 5046 9818
rect 5046 9766 5052 9818
rect 5076 9766 5098 9818
rect 5098 9766 5110 9818
rect 5110 9766 5132 9818
rect 5156 9766 5162 9818
rect 5162 9766 5174 9818
rect 5174 9766 5212 9818
rect 5236 9766 5238 9818
rect 5238 9766 5290 9818
rect 5290 9766 5292 9818
rect 4916 9764 4972 9766
rect 4996 9764 5052 9766
rect 5076 9764 5132 9766
rect 5156 9764 5212 9766
rect 5236 9764 5292 9766
rect 6182 13388 6238 13424
rect 6182 13368 6184 13388
rect 6184 13368 6236 13388
rect 6236 13368 6238 13388
rect 7194 13368 7250 13424
rect 4916 8730 4972 8732
rect 4996 8730 5052 8732
rect 5076 8730 5132 8732
rect 5156 8730 5212 8732
rect 5236 8730 5292 8732
rect 4916 8678 4918 8730
rect 4918 8678 4970 8730
rect 4970 8678 4972 8730
rect 4996 8678 5034 8730
rect 5034 8678 5046 8730
rect 5046 8678 5052 8730
rect 5076 8678 5098 8730
rect 5098 8678 5110 8730
rect 5110 8678 5132 8730
rect 5156 8678 5162 8730
rect 5162 8678 5174 8730
rect 5174 8678 5212 8730
rect 5236 8678 5238 8730
rect 5238 8678 5290 8730
rect 5290 8678 5292 8730
rect 4916 8676 4972 8678
rect 4996 8676 5052 8678
rect 5076 8676 5132 8678
rect 5156 8676 5212 8678
rect 5236 8676 5292 8678
rect 5998 11772 6000 11792
rect 6000 11772 6052 11792
rect 6052 11772 6054 11792
rect 5998 11736 6054 11772
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 6090 10920 6146 10976
rect 4986 7828 4988 7848
rect 4988 7828 5040 7848
rect 5040 7828 5042 7848
rect 4986 7792 5042 7828
rect 4916 7642 4972 7644
rect 4996 7642 5052 7644
rect 5076 7642 5132 7644
rect 5156 7642 5212 7644
rect 5236 7642 5292 7644
rect 4916 7590 4918 7642
rect 4918 7590 4970 7642
rect 4970 7590 4972 7642
rect 4996 7590 5034 7642
rect 5034 7590 5046 7642
rect 5046 7590 5052 7642
rect 5076 7590 5098 7642
rect 5098 7590 5110 7642
rect 5110 7590 5132 7642
rect 5156 7590 5162 7642
rect 5162 7590 5174 7642
rect 5174 7590 5212 7642
rect 5236 7590 5238 7642
rect 5238 7590 5290 7642
rect 5290 7590 5292 7642
rect 4916 7588 4972 7590
rect 4996 7588 5052 7590
rect 5076 7588 5132 7590
rect 5156 7588 5212 7590
rect 5236 7588 5292 7590
rect 4916 6554 4972 6556
rect 4996 6554 5052 6556
rect 5076 6554 5132 6556
rect 5156 6554 5212 6556
rect 5236 6554 5292 6556
rect 4916 6502 4918 6554
rect 4918 6502 4970 6554
rect 4970 6502 4972 6554
rect 4996 6502 5034 6554
rect 5034 6502 5046 6554
rect 5046 6502 5052 6554
rect 5076 6502 5098 6554
rect 5098 6502 5110 6554
rect 5110 6502 5132 6554
rect 5156 6502 5162 6554
rect 5162 6502 5174 6554
rect 5174 6502 5212 6554
rect 5236 6502 5238 6554
rect 5238 6502 5290 6554
rect 5290 6502 5292 6554
rect 4916 6500 4972 6502
rect 4996 6500 5052 6502
rect 5076 6500 5132 6502
rect 5156 6500 5212 6502
rect 5236 6500 5292 6502
rect 4916 5466 4972 5468
rect 4996 5466 5052 5468
rect 5076 5466 5132 5468
rect 5156 5466 5212 5468
rect 5236 5466 5292 5468
rect 4916 5414 4918 5466
rect 4918 5414 4970 5466
rect 4970 5414 4972 5466
rect 4996 5414 5034 5466
rect 5034 5414 5046 5466
rect 5046 5414 5052 5466
rect 5076 5414 5098 5466
rect 5098 5414 5110 5466
rect 5110 5414 5132 5466
rect 5156 5414 5162 5466
rect 5162 5414 5174 5466
rect 5174 5414 5212 5466
rect 5236 5414 5238 5466
rect 5238 5414 5290 5466
rect 5290 5414 5292 5466
rect 4916 5412 4972 5414
rect 4996 5412 5052 5414
rect 5076 5412 5132 5414
rect 5156 5412 5212 5414
rect 5236 5412 5292 5414
rect 4434 4276 4490 4312
rect 4434 4256 4436 4276
rect 4436 4256 4488 4276
rect 4488 4256 4490 4276
rect 4434 3984 4490 4040
rect 4916 4378 4972 4380
rect 4996 4378 5052 4380
rect 5076 4378 5132 4380
rect 5156 4378 5212 4380
rect 5236 4378 5292 4380
rect 4916 4326 4918 4378
rect 4918 4326 4970 4378
rect 4970 4326 4972 4378
rect 4996 4326 5034 4378
rect 5034 4326 5046 4378
rect 5046 4326 5052 4378
rect 5076 4326 5098 4378
rect 5098 4326 5110 4378
rect 5110 4326 5132 4378
rect 5156 4326 5162 4378
rect 5162 4326 5174 4378
rect 5174 4326 5212 4378
rect 5236 4326 5238 4378
rect 5238 4326 5290 4378
rect 5290 4326 5292 4378
rect 4916 4324 4972 4326
rect 4996 4324 5052 4326
rect 5076 4324 5132 4326
rect 5156 4324 5212 4326
rect 5236 4324 5292 4326
rect 6918 11192 6974 11248
rect 6826 10784 6882 10840
rect 6826 10668 6882 10704
rect 6826 10648 6828 10668
rect 6828 10648 6880 10668
rect 6880 10648 6882 10668
rect 7654 11600 7710 11656
rect 7194 10920 7250 10976
rect 7378 10648 7434 10704
rect 6918 6740 6920 6760
rect 6920 6740 6972 6760
rect 6972 6740 6974 6760
rect 6918 6704 6974 6740
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 7930 11192 7986 11248
rect 10916 14170 10972 14172
rect 10996 14170 11052 14172
rect 11076 14170 11132 14172
rect 11156 14170 11212 14172
rect 11236 14170 11292 14172
rect 10916 14118 10918 14170
rect 10918 14118 10970 14170
rect 10970 14118 10972 14170
rect 10996 14118 11034 14170
rect 11034 14118 11046 14170
rect 11046 14118 11052 14170
rect 11076 14118 11098 14170
rect 11098 14118 11110 14170
rect 11110 14118 11132 14170
rect 11156 14118 11162 14170
rect 11162 14118 11174 14170
rect 11174 14118 11212 14170
rect 11236 14118 11238 14170
rect 11238 14118 11290 14170
rect 11290 14118 11292 14170
rect 10916 14116 10972 14118
rect 10996 14116 11052 14118
rect 11076 14116 11132 14118
rect 11156 14116 11212 14118
rect 11236 14116 11292 14118
rect 10138 13776 10194 13832
rect 10046 13640 10102 13696
rect 7930 10784 7986 10840
rect 8022 10648 8078 10704
rect 8482 11056 8538 11112
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 9034 10784 9090 10840
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 4916 3290 4972 3292
rect 4996 3290 5052 3292
rect 5076 3290 5132 3292
rect 5156 3290 5212 3292
rect 5236 3290 5292 3292
rect 4916 3238 4918 3290
rect 4918 3238 4970 3290
rect 4970 3238 4972 3290
rect 4996 3238 5034 3290
rect 5034 3238 5046 3290
rect 5046 3238 5052 3290
rect 5076 3238 5098 3290
rect 5098 3238 5110 3290
rect 5110 3238 5132 3290
rect 5156 3238 5162 3290
rect 5162 3238 5174 3290
rect 5174 3238 5212 3290
rect 5236 3238 5238 3290
rect 5238 3238 5290 3290
rect 5290 3238 5292 3290
rect 4916 3236 4972 3238
rect 4996 3236 5052 3238
rect 5076 3236 5132 3238
rect 5156 3236 5212 3238
rect 5236 3236 5292 3238
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 10322 12280 10378 12336
rect 9678 10376 9734 10432
rect 9310 8336 9366 8392
rect 9678 9580 9734 9616
rect 9678 9560 9680 9580
rect 9680 9560 9732 9580
rect 9732 9560 9734 9580
rect 9954 11192 10010 11248
rect 9862 9424 9918 9480
rect 9770 9152 9826 9208
rect 9770 9036 9826 9072
rect 9770 9016 9772 9036
rect 9772 9016 9824 9036
rect 9824 9016 9826 9036
rect 8666 7792 8722 7848
rect 10230 12144 10286 12200
rect 10046 10104 10102 10160
rect 10916 13082 10972 13084
rect 10996 13082 11052 13084
rect 11076 13082 11132 13084
rect 11156 13082 11212 13084
rect 11236 13082 11292 13084
rect 10916 13030 10918 13082
rect 10918 13030 10970 13082
rect 10970 13030 10972 13082
rect 10996 13030 11034 13082
rect 11034 13030 11046 13082
rect 11046 13030 11052 13082
rect 11076 13030 11098 13082
rect 11098 13030 11110 13082
rect 11110 13030 11132 13082
rect 11156 13030 11162 13082
rect 11162 13030 11174 13082
rect 11174 13030 11212 13082
rect 11236 13030 11238 13082
rect 11238 13030 11290 13082
rect 11290 13030 11292 13082
rect 10916 13028 10972 13030
rect 10996 13028 11052 13030
rect 11076 13028 11132 13030
rect 11156 13028 11212 13030
rect 11236 13028 11292 13030
rect 10874 12280 10930 12336
rect 10966 12144 11022 12200
rect 10916 11994 10972 11996
rect 10996 11994 11052 11996
rect 11076 11994 11132 11996
rect 11156 11994 11212 11996
rect 11236 11994 11292 11996
rect 10916 11942 10918 11994
rect 10918 11942 10970 11994
rect 10970 11942 10972 11994
rect 10996 11942 11034 11994
rect 11034 11942 11046 11994
rect 11046 11942 11052 11994
rect 11076 11942 11098 11994
rect 11098 11942 11110 11994
rect 11110 11942 11132 11994
rect 11156 11942 11162 11994
rect 11162 11942 11174 11994
rect 11174 11942 11212 11994
rect 11236 11942 11238 11994
rect 11238 11942 11290 11994
rect 11290 11942 11292 11994
rect 10916 11940 10972 11942
rect 10996 11940 11052 11942
rect 11076 11940 11132 11942
rect 11156 11940 11212 11942
rect 11236 11940 11292 11942
rect 11242 11464 11298 11520
rect 11150 11328 11206 11384
rect 11426 11192 11482 11248
rect 10782 11056 10838 11112
rect 10916 10906 10972 10908
rect 10996 10906 11052 10908
rect 11076 10906 11132 10908
rect 11156 10906 11212 10908
rect 11236 10906 11292 10908
rect 10916 10854 10918 10906
rect 10918 10854 10970 10906
rect 10970 10854 10972 10906
rect 10996 10854 11034 10906
rect 11034 10854 11046 10906
rect 11046 10854 11052 10906
rect 11076 10854 11098 10906
rect 11098 10854 11110 10906
rect 11110 10854 11132 10906
rect 11156 10854 11162 10906
rect 11162 10854 11174 10906
rect 11174 10854 11212 10906
rect 11236 10854 11238 10906
rect 11238 10854 11290 10906
rect 11290 10854 11292 10906
rect 10916 10852 10972 10854
rect 10996 10852 11052 10854
rect 11076 10852 11132 10854
rect 11156 10852 11212 10854
rect 11236 10852 11292 10854
rect 10690 10512 10746 10568
rect 11058 10512 11114 10568
rect 10598 10376 10654 10432
rect 10782 10376 10838 10432
rect 10506 9288 10562 9344
rect 10230 8880 10286 8936
rect 10690 10104 10746 10160
rect 11334 10512 11390 10568
rect 10916 9818 10972 9820
rect 10996 9818 11052 9820
rect 11076 9818 11132 9820
rect 11156 9818 11212 9820
rect 11236 9818 11292 9820
rect 10916 9766 10918 9818
rect 10918 9766 10970 9818
rect 10970 9766 10972 9818
rect 10996 9766 11034 9818
rect 11034 9766 11046 9818
rect 11046 9766 11052 9818
rect 11076 9766 11098 9818
rect 11098 9766 11110 9818
rect 11110 9766 11132 9818
rect 11156 9766 11162 9818
rect 11162 9766 11174 9818
rect 11174 9766 11212 9818
rect 11236 9766 11238 9818
rect 11238 9766 11290 9818
rect 11290 9766 11292 9818
rect 10916 9764 10972 9766
rect 10996 9764 11052 9766
rect 11076 9764 11132 9766
rect 11156 9764 11212 9766
rect 11236 9764 11292 9766
rect 10690 9152 10746 9208
rect 10598 8744 10654 8800
rect 9402 6704 9458 6760
rect 9954 7928 10010 7984
rect 9678 6296 9734 6352
rect 9770 5752 9826 5808
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 11058 9052 11060 9072
rect 11060 9052 11112 9072
rect 11112 9052 11114 9072
rect 11058 9016 11114 9052
rect 11334 8880 11390 8936
rect 10916 8730 10972 8732
rect 10996 8730 11052 8732
rect 11076 8730 11132 8732
rect 11156 8730 11212 8732
rect 11236 8730 11292 8732
rect 10916 8678 10918 8730
rect 10918 8678 10970 8730
rect 10970 8678 10972 8730
rect 10996 8678 11034 8730
rect 11034 8678 11046 8730
rect 11046 8678 11052 8730
rect 11076 8678 11098 8730
rect 11098 8678 11110 8730
rect 11110 8678 11132 8730
rect 11156 8678 11162 8730
rect 11162 8678 11174 8730
rect 11174 8678 11212 8730
rect 11236 8678 11238 8730
rect 11238 8678 11290 8730
rect 11290 8678 11292 8730
rect 10916 8676 10972 8678
rect 10996 8676 11052 8678
rect 11076 8676 11132 8678
rect 11156 8676 11212 8678
rect 11236 8676 11292 8678
rect 11150 8492 11206 8528
rect 11150 8472 11152 8492
rect 11152 8472 11204 8492
rect 11204 8472 11206 8492
rect 10916 7642 10972 7644
rect 10996 7642 11052 7644
rect 11076 7642 11132 7644
rect 11156 7642 11212 7644
rect 11236 7642 11292 7644
rect 10916 7590 10918 7642
rect 10918 7590 10970 7642
rect 10970 7590 10972 7642
rect 10996 7590 11034 7642
rect 11034 7590 11046 7642
rect 11046 7590 11052 7642
rect 11076 7590 11098 7642
rect 11098 7590 11110 7642
rect 11110 7590 11132 7642
rect 11156 7590 11162 7642
rect 11162 7590 11174 7642
rect 11174 7590 11212 7642
rect 11236 7590 11238 7642
rect 11238 7590 11290 7642
rect 11290 7590 11292 7642
rect 10916 7588 10972 7590
rect 10996 7588 11052 7590
rect 11076 7588 11132 7590
rect 11156 7588 11212 7590
rect 11236 7588 11292 7590
rect 11794 10512 11850 10568
rect 12162 12144 12218 12200
rect 11610 9424 11666 9480
rect 11610 9152 11666 9208
rect 10046 6160 10102 6216
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 10916 6554 10972 6556
rect 10996 6554 11052 6556
rect 11076 6554 11132 6556
rect 11156 6554 11212 6556
rect 11236 6554 11292 6556
rect 10916 6502 10918 6554
rect 10918 6502 10970 6554
rect 10970 6502 10972 6554
rect 10996 6502 11034 6554
rect 11034 6502 11046 6554
rect 11046 6502 11052 6554
rect 11076 6502 11098 6554
rect 11098 6502 11110 6554
rect 11110 6502 11132 6554
rect 11156 6502 11162 6554
rect 11162 6502 11174 6554
rect 11174 6502 11212 6554
rect 11236 6502 11238 6554
rect 11238 6502 11290 6554
rect 11290 6502 11292 6554
rect 10916 6500 10972 6502
rect 10996 6500 11052 6502
rect 11076 6500 11132 6502
rect 11156 6500 11212 6502
rect 11236 6500 11292 6502
rect 10916 5466 10972 5468
rect 10996 5466 11052 5468
rect 11076 5466 11132 5468
rect 11156 5466 11212 5468
rect 11236 5466 11292 5468
rect 10916 5414 10918 5466
rect 10918 5414 10970 5466
rect 10970 5414 10972 5466
rect 10996 5414 11034 5466
rect 11034 5414 11046 5466
rect 11046 5414 11052 5466
rect 11076 5414 11098 5466
rect 11098 5414 11110 5466
rect 11110 5414 11132 5466
rect 11156 5414 11162 5466
rect 11162 5414 11174 5466
rect 11174 5414 11212 5466
rect 11236 5414 11238 5466
rect 11238 5414 11290 5466
rect 11290 5414 11292 5466
rect 10916 5412 10972 5414
rect 10996 5412 11052 5414
rect 11076 5412 11132 5414
rect 11156 5412 11212 5414
rect 11236 5412 11292 5414
rect 12162 11756 12218 11792
rect 12162 11736 12164 11756
rect 12164 11736 12216 11756
rect 12216 11736 12218 11756
rect 12530 11464 12586 11520
rect 12714 11328 12770 11384
rect 12346 11092 12348 11112
rect 12348 11092 12400 11112
rect 12400 11092 12402 11112
rect 12346 11056 12402 11092
rect 12070 10376 12126 10432
rect 12070 5788 12072 5808
rect 12072 5788 12124 5808
rect 12124 5788 12126 5808
rect 12070 5752 12126 5788
rect 10916 4378 10972 4380
rect 10996 4378 11052 4380
rect 11076 4378 11132 4380
rect 11156 4378 11212 4380
rect 11236 4378 11292 4380
rect 10916 4326 10918 4378
rect 10918 4326 10970 4378
rect 10970 4326 10972 4378
rect 10996 4326 11034 4378
rect 11034 4326 11046 4378
rect 11046 4326 11052 4378
rect 11076 4326 11098 4378
rect 11098 4326 11110 4378
rect 11110 4326 11132 4378
rect 11156 4326 11162 4378
rect 11162 4326 11174 4378
rect 11174 4326 11212 4378
rect 11236 4326 11238 4378
rect 11238 4326 11290 4378
rect 11290 4326 11292 4378
rect 10916 4324 10972 4326
rect 10996 4324 11052 4326
rect 11076 4324 11132 4326
rect 11156 4324 11212 4326
rect 11236 4324 11292 4326
rect 10138 3984 10194 4040
rect 4916 2202 4972 2204
rect 4996 2202 5052 2204
rect 5076 2202 5132 2204
rect 5156 2202 5212 2204
rect 5236 2202 5292 2204
rect 4916 2150 4918 2202
rect 4918 2150 4970 2202
rect 4970 2150 4972 2202
rect 4996 2150 5034 2202
rect 5034 2150 5046 2202
rect 5046 2150 5052 2202
rect 5076 2150 5098 2202
rect 5098 2150 5110 2202
rect 5110 2150 5132 2202
rect 5156 2150 5162 2202
rect 5162 2150 5174 2202
rect 5174 2150 5212 2202
rect 5236 2150 5238 2202
rect 5238 2150 5290 2202
rect 5290 2150 5292 2202
rect 4916 2148 4972 2150
rect 4996 2148 5052 2150
rect 5076 2148 5132 2150
rect 5156 2148 5212 2150
rect 5236 2148 5292 2150
rect 10916 3290 10972 3292
rect 10996 3290 11052 3292
rect 11076 3290 11132 3292
rect 11156 3290 11212 3292
rect 11236 3290 11292 3292
rect 10916 3238 10918 3290
rect 10918 3238 10970 3290
rect 10970 3238 10972 3290
rect 10996 3238 11034 3290
rect 11034 3238 11046 3290
rect 11046 3238 11052 3290
rect 11076 3238 11098 3290
rect 11098 3238 11110 3290
rect 11110 3238 11132 3290
rect 11156 3238 11162 3290
rect 11162 3238 11174 3290
rect 11174 3238 11212 3290
rect 11236 3238 11238 3290
rect 11238 3238 11290 3290
rect 11290 3238 11292 3290
rect 10916 3236 10972 3238
rect 10996 3236 11052 3238
rect 11076 3236 11132 3238
rect 11156 3236 11212 3238
rect 11236 3236 11292 3238
rect 10916 2202 10972 2204
rect 10996 2202 11052 2204
rect 11076 2202 11132 2204
rect 11156 2202 11212 2204
rect 11236 2202 11292 2204
rect 10916 2150 10918 2202
rect 10918 2150 10970 2202
rect 10970 2150 10972 2202
rect 10996 2150 11034 2202
rect 11034 2150 11046 2202
rect 11046 2150 11052 2202
rect 11076 2150 11098 2202
rect 11098 2150 11110 2202
rect 11110 2150 11132 2202
rect 11156 2150 11162 2202
rect 11162 2150 11174 2202
rect 11174 2150 11212 2202
rect 11236 2150 11238 2202
rect 11238 2150 11290 2202
rect 11290 2150 11292 2202
rect 10916 2148 10972 2150
rect 10996 2148 11052 2150
rect 11076 2148 11132 2150
rect 11156 2148 11212 2150
rect 11236 2148 11292 2150
<< metal3 >>
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 4906 14176 5302 14177
rect 4906 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5302 14176
rect 4906 14111 5302 14112
rect 10906 14176 11302 14177
rect 10906 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11302 14176
rect 10906 14111 11302 14112
rect 9990 13772 9996 13836
rect 10060 13834 10066 13836
rect 10133 13834 10199 13837
rect 10060 13832 10199 13834
rect 10060 13776 10138 13832
rect 10194 13776 10199 13832
rect 10060 13774 10199 13776
rect 10060 13772 10066 13774
rect 10133 13771 10199 13774
rect 10041 13698 10107 13701
rect 10174 13698 10180 13700
rect 10041 13696 10180 13698
rect 10041 13640 10046 13696
rect 10102 13640 10180 13696
rect 10041 13638 10180 13640
rect 10041 13635 10107 13638
rect 10174 13636 10180 13638
rect 10244 13636 10250 13700
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 3417 13426 3483 13429
rect 4429 13426 4495 13429
rect 3417 13424 4495 13426
rect 3417 13368 3422 13424
rect 3478 13368 4434 13424
rect 4490 13368 4495 13424
rect 3417 13366 4495 13368
rect 3417 13363 3483 13366
rect 4429 13363 4495 13366
rect 6177 13426 6243 13429
rect 7189 13426 7255 13429
rect 6177 13424 7255 13426
rect 6177 13368 6182 13424
rect 6238 13368 7194 13424
rect 7250 13368 7255 13424
rect 6177 13366 7255 13368
rect 6177 13363 6243 13366
rect 7189 13363 7255 13366
rect 4906 13088 5302 13089
rect 4906 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5302 13088
rect 4906 13023 5302 13024
rect 10906 13088 11302 13089
rect 10906 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11302 13088
rect 10906 13023 11302 13024
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 10317 12338 10383 12341
rect 10869 12338 10935 12341
rect 10317 12336 10935 12338
rect 10317 12280 10322 12336
rect 10378 12280 10874 12336
rect 10930 12280 10935 12336
rect 10317 12278 10935 12280
rect 10317 12275 10383 12278
rect 10869 12275 10935 12278
rect 10225 12202 10291 12205
rect 10961 12202 11027 12205
rect 12157 12202 12223 12205
rect 10225 12200 12223 12202
rect 10225 12144 10230 12200
rect 10286 12144 10966 12200
rect 11022 12144 12162 12200
rect 12218 12144 12223 12200
rect 10225 12142 12223 12144
rect 10225 12139 10291 12142
rect 10961 12139 11027 12142
rect 12157 12139 12223 12142
rect 4906 12000 5302 12001
rect 4906 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5302 12000
rect 4906 11935 5302 11936
rect 10906 12000 11302 12001
rect 10906 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11302 12000
rect 10906 11935 11302 11936
rect 4429 11794 4495 11797
rect 5993 11794 6059 11797
rect 4429 11792 6059 11794
rect 4429 11736 4434 11792
rect 4490 11736 5998 11792
rect 6054 11736 6059 11792
rect 4429 11734 6059 11736
rect 4429 11731 4495 11734
rect 5993 11731 6059 11734
rect 9990 11732 9996 11796
rect 10060 11794 10066 11796
rect 12157 11794 12223 11797
rect 10060 11792 12223 11794
rect 10060 11736 12162 11792
rect 12218 11736 12223 11792
rect 10060 11734 12223 11736
rect 10060 11732 10066 11734
rect 12157 11731 12223 11734
rect 5073 11658 5139 11661
rect 7649 11658 7715 11661
rect 5073 11656 7715 11658
rect 5073 11600 5078 11656
rect 5134 11600 7654 11656
rect 7710 11600 7715 11656
rect 5073 11598 7715 11600
rect 5073 11595 5139 11598
rect 7649 11595 7715 11598
rect 4245 11524 4311 11525
rect 4245 11522 4292 11524
rect 4200 11520 4292 11522
rect 4200 11464 4250 11520
rect 4200 11462 4292 11464
rect 4245 11460 4292 11462
rect 4356 11460 4362 11524
rect 11237 11522 11303 11525
rect 12525 11522 12591 11525
rect 11237 11520 12591 11522
rect 11237 11464 11242 11520
rect 11298 11464 12530 11520
rect 12586 11464 12591 11520
rect 11237 11462 12591 11464
rect 4245 11459 4311 11460
rect 11237 11459 11303 11462
rect 12525 11459 12591 11462
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 4981 11386 5047 11389
rect 5349 11386 5415 11389
rect 4981 11384 5415 11386
rect 4981 11328 4986 11384
rect 5042 11328 5354 11384
rect 5410 11328 5415 11384
rect 4981 11326 5415 11328
rect 4981 11323 5047 11326
rect 5349 11323 5415 11326
rect 11145 11386 11211 11389
rect 12709 11386 12775 11389
rect 11145 11384 12775 11386
rect 11145 11328 11150 11384
rect 11206 11328 12714 11384
rect 12770 11328 12775 11384
rect 11145 11326 12775 11328
rect 11145 11323 11211 11326
rect 12709 11323 12775 11326
rect 6913 11250 6979 11253
rect 7925 11250 7991 11253
rect 6913 11248 7991 11250
rect 6913 11192 6918 11248
rect 6974 11192 7930 11248
rect 7986 11192 7991 11248
rect 6913 11190 7991 11192
rect 6913 11187 6979 11190
rect 7925 11187 7991 11190
rect 9949 11250 10015 11253
rect 11421 11250 11487 11253
rect 9949 11248 11487 11250
rect 9949 11192 9954 11248
rect 10010 11192 11426 11248
rect 11482 11192 11487 11248
rect 9949 11190 11487 11192
rect 9949 11187 10015 11190
rect 11421 11187 11487 11190
rect 4981 11114 5047 11117
rect 8477 11114 8543 11117
rect 4981 11112 8543 11114
rect 4981 11056 4986 11112
rect 5042 11056 8482 11112
rect 8538 11056 8543 11112
rect 4981 11054 8543 11056
rect 4981 11051 5047 11054
rect 8477 11051 8543 11054
rect 10777 11114 10843 11117
rect 12341 11114 12407 11117
rect 10777 11112 12407 11114
rect 10777 11056 10782 11112
rect 10838 11056 12346 11112
rect 12402 11056 12407 11112
rect 10777 11054 12407 11056
rect 10777 11051 10843 11054
rect 12341 11051 12407 11054
rect 6085 10978 6151 10981
rect 7189 10978 7255 10981
rect 6085 10976 7255 10978
rect 6085 10920 6090 10976
rect 6146 10920 7194 10976
rect 7250 10920 7255 10976
rect 6085 10918 7255 10920
rect 6085 10915 6151 10918
rect 7189 10915 7255 10918
rect 4906 10912 5302 10913
rect 4906 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5302 10912
rect 4906 10847 5302 10848
rect 10906 10912 11302 10913
rect 10906 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11302 10912
rect 10906 10847 11302 10848
rect 6821 10842 6887 10845
rect 7925 10842 7991 10845
rect 9029 10842 9095 10845
rect 6821 10840 9095 10842
rect 6821 10784 6826 10840
rect 6882 10784 7930 10840
rect 7986 10784 9034 10840
rect 9090 10784 9095 10840
rect 6821 10782 9095 10784
rect 6821 10779 6887 10782
rect 7925 10779 7991 10782
rect 9029 10779 9095 10782
rect 6821 10706 6887 10709
rect 7373 10706 7439 10709
rect 8017 10706 8083 10709
rect 6821 10704 8083 10706
rect 6821 10648 6826 10704
rect 6882 10648 7378 10704
rect 7434 10648 8022 10704
rect 8078 10648 8083 10704
rect 6821 10646 8083 10648
rect 6821 10643 6887 10646
rect 7373 10643 7439 10646
rect 8017 10643 8083 10646
rect 10685 10570 10751 10573
rect 11053 10570 11119 10573
rect 10685 10568 11119 10570
rect 10685 10512 10690 10568
rect 10746 10512 11058 10568
rect 11114 10512 11119 10568
rect 10685 10510 11119 10512
rect 10685 10507 10751 10510
rect 11053 10507 11119 10510
rect 11329 10570 11395 10573
rect 11789 10570 11855 10573
rect 11329 10568 11855 10570
rect 11329 10512 11334 10568
rect 11390 10512 11794 10568
rect 11850 10512 11855 10568
rect 11329 10510 11855 10512
rect 11329 10507 11395 10510
rect 11789 10507 11855 10510
rect 9673 10434 9739 10437
rect 10593 10434 10659 10437
rect 9673 10432 10659 10434
rect 9673 10376 9678 10432
rect 9734 10376 10598 10432
rect 10654 10376 10659 10432
rect 9673 10374 10659 10376
rect 9673 10371 9739 10374
rect 10593 10371 10659 10374
rect 10777 10434 10843 10437
rect 12065 10434 12131 10437
rect 10777 10432 12131 10434
rect 10777 10376 10782 10432
rect 10838 10376 12070 10432
rect 12126 10376 12131 10432
rect 10777 10374 12131 10376
rect 10777 10371 10843 10374
rect 12065 10371 12131 10374
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 10041 10162 10107 10165
rect 10685 10162 10751 10165
rect 10041 10160 10751 10162
rect 10041 10104 10046 10160
rect 10102 10104 10690 10160
rect 10746 10104 10751 10160
rect 10041 10102 10751 10104
rect 10041 10099 10107 10102
rect 10685 10099 10751 10102
rect 4906 9824 5302 9825
rect 4906 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5302 9824
rect 4906 9759 5302 9760
rect 10906 9824 11302 9825
rect 10906 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11302 9824
rect 10906 9759 11302 9760
rect 9673 9618 9739 9621
rect 9630 9616 9739 9618
rect 9630 9560 9678 9616
rect 9734 9560 9739 9616
rect 9630 9555 9739 9560
rect 9630 9346 9690 9555
rect 9857 9482 9923 9485
rect 11605 9482 11671 9485
rect 9857 9480 11671 9482
rect 9857 9424 9862 9480
rect 9918 9424 11610 9480
rect 11666 9424 11671 9480
rect 9857 9422 11671 9424
rect 9857 9419 9923 9422
rect 11605 9419 11671 9422
rect 10501 9346 10567 9349
rect 9630 9344 10567 9346
rect 9630 9288 10506 9344
rect 10562 9288 10567 9344
rect 9630 9286 10567 9288
rect 10501 9283 10567 9286
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 9765 9210 9831 9213
rect 10685 9210 10751 9213
rect 11605 9210 11671 9213
rect 9765 9208 11671 9210
rect 9765 9152 9770 9208
rect 9826 9152 10690 9208
rect 10746 9152 11610 9208
rect 11666 9152 11671 9208
rect 9765 9150 11671 9152
rect 9765 9147 9831 9150
rect 10685 9147 10751 9150
rect 11605 9147 11671 9150
rect 9765 9074 9831 9077
rect 11053 9074 11119 9077
rect 9765 9072 11119 9074
rect 9765 9016 9770 9072
rect 9826 9016 11058 9072
rect 11114 9016 11119 9072
rect 9765 9014 11119 9016
rect 9765 9011 9831 9014
rect 11053 9011 11119 9014
rect 10225 8938 10291 8941
rect 11329 8938 11395 8941
rect 10225 8936 11395 8938
rect 10225 8880 10230 8936
rect 10286 8880 11334 8936
rect 11390 8880 11395 8936
rect 10225 8878 11395 8880
rect 10225 8875 10291 8878
rect 11329 8875 11395 8878
rect 10593 8802 10659 8805
rect 10593 8800 10794 8802
rect 10593 8744 10598 8800
rect 10654 8744 10794 8800
rect 10593 8742 10794 8744
rect 10593 8739 10659 8742
rect 4906 8736 5302 8737
rect 4906 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5302 8736
rect 4906 8671 5302 8672
rect 10734 8530 10794 8742
rect 10906 8736 11302 8737
rect 10906 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11302 8736
rect 10906 8671 11302 8672
rect 11145 8530 11211 8533
rect 10734 8528 11211 8530
rect 10734 8472 11150 8528
rect 11206 8472 11211 8528
rect 10734 8470 11211 8472
rect 11145 8467 11211 8470
rect 2129 8394 2195 8397
rect 9305 8394 9371 8397
rect 2129 8392 9371 8394
rect 2129 8336 2134 8392
rect 2190 8336 9310 8392
rect 9366 8336 9371 8392
rect 2129 8334 9371 8336
rect 2129 8331 2195 8334
rect 9305 8331 9371 8334
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 9949 7988 10015 7989
rect 9949 7986 9996 7988
rect 9904 7984 9996 7986
rect 9904 7928 9954 7984
rect 9904 7926 9996 7928
rect 9949 7924 9996 7926
rect 10060 7924 10066 7988
rect 9949 7923 10015 7924
rect 4981 7850 5047 7853
rect 8661 7850 8727 7853
rect 4981 7848 8727 7850
rect 4981 7792 4986 7848
rect 5042 7792 8666 7848
rect 8722 7792 8727 7848
rect 4981 7790 8727 7792
rect 4981 7787 5047 7790
rect 8661 7787 8727 7790
rect 4906 7648 5302 7649
rect 4906 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5302 7648
rect 4906 7583 5302 7584
rect 10906 7648 11302 7649
rect 10906 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11302 7648
rect 10906 7583 11302 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 6913 6762 6979 6765
rect 9397 6762 9463 6765
rect 6913 6760 9463 6762
rect 6913 6704 6918 6760
rect 6974 6704 9402 6760
rect 9458 6704 9463 6760
rect 6913 6702 9463 6704
rect 6913 6699 6979 6702
rect 9397 6699 9463 6702
rect 4906 6560 5302 6561
rect 4906 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5302 6560
rect 4906 6495 5302 6496
rect 10906 6560 11302 6561
rect 10906 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11302 6560
rect 10906 6495 11302 6496
rect 9673 6354 9739 6357
rect 9673 6352 10058 6354
rect 9673 6296 9678 6352
rect 9734 6296 10058 6352
rect 9673 6294 10058 6296
rect 9673 6291 9739 6294
rect 9998 6221 10058 6294
rect 9998 6216 10107 6221
rect 9998 6160 10046 6216
rect 10102 6160 10107 6216
rect 9998 6158 10107 6160
rect 10041 6155 10107 6158
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 9765 5810 9831 5813
rect 12065 5810 12131 5813
rect 9765 5808 12131 5810
rect 9765 5752 9770 5808
rect 9826 5752 12070 5808
rect 12126 5752 12131 5808
rect 9765 5750 12131 5752
rect 9765 5747 9831 5750
rect 12065 5747 12131 5750
rect 4906 5472 5302 5473
rect 4906 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5302 5472
rect 4906 5407 5302 5408
rect 10906 5472 11302 5473
rect 10906 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11302 5472
rect 10906 5407 11302 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 4906 4384 5302 4385
rect 4906 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5302 4384
rect 4906 4319 5302 4320
rect 10906 4384 11302 4385
rect 10906 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11302 4384
rect 10906 4319 11302 4320
rect 3969 4314 4035 4317
rect 4429 4314 4495 4317
rect 3969 4312 4495 4314
rect 3969 4256 3974 4312
rect 4030 4256 4434 4312
rect 4490 4256 4495 4312
rect 3969 4254 4495 4256
rect 3969 4251 4035 4254
rect 4429 4251 4495 4254
rect 4286 3980 4292 4044
rect 4356 4042 4362 4044
rect 4429 4042 4495 4045
rect 10133 4044 10199 4045
rect 10133 4042 10180 4044
rect 4356 4040 4495 4042
rect 4356 3984 4434 4040
rect 4490 3984 4495 4040
rect 4356 3982 4495 3984
rect 10088 4040 10180 4042
rect 10088 3984 10138 4040
rect 10088 3982 10180 3984
rect 4356 3980 4362 3982
rect 4429 3979 4495 3982
rect 10133 3980 10180 3982
rect 10244 3980 10250 4044
rect 10133 3979 10199 3980
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 4906 3296 5302 3297
rect 4906 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5302 3296
rect 4906 3231 5302 3232
rect 10906 3296 11302 3297
rect 10906 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11302 3296
rect 10906 3231 11302 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 4906 2208 5302 2209
rect 4906 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5302 2208
rect 4906 2143 5302 2144
rect 10906 2208 11302 2209
rect 10906 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11302 2208
rect 10906 2143 11302 2144
<< via3 >>
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 4912 14172 4976 14176
rect 4912 14116 4916 14172
rect 4916 14116 4972 14172
rect 4972 14116 4976 14172
rect 4912 14112 4976 14116
rect 4992 14172 5056 14176
rect 4992 14116 4996 14172
rect 4996 14116 5052 14172
rect 5052 14116 5056 14172
rect 4992 14112 5056 14116
rect 5072 14172 5136 14176
rect 5072 14116 5076 14172
rect 5076 14116 5132 14172
rect 5132 14116 5136 14172
rect 5072 14112 5136 14116
rect 5152 14172 5216 14176
rect 5152 14116 5156 14172
rect 5156 14116 5212 14172
rect 5212 14116 5216 14172
rect 5152 14112 5216 14116
rect 5232 14172 5296 14176
rect 5232 14116 5236 14172
rect 5236 14116 5292 14172
rect 5292 14116 5296 14172
rect 5232 14112 5296 14116
rect 10912 14172 10976 14176
rect 10912 14116 10916 14172
rect 10916 14116 10972 14172
rect 10972 14116 10976 14172
rect 10912 14112 10976 14116
rect 10992 14172 11056 14176
rect 10992 14116 10996 14172
rect 10996 14116 11052 14172
rect 11052 14116 11056 14172
rect 10992 14112 11056 14116
rect 11072 14172 11136 14176
rect 11072 14116 11076 14172
rect 11076 14116 11132 14172
rect 11132 14116 11136 14172
rect 11072 14112 11136 14116
rect 11152 14172 11216 14176
rect 11152 14116 11156 14172
rect 11156 14116 11212 14172
rect 11212 14116 11216 14172
rect 11152 14112 11216 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 9996 13772 10060 13836
rect 10180 13636 10244 13700
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 4912 13084 4976 13088
rect 4912 13028 4916 13084
rect 4916 13028 4972 13084
rect 4972 13028 4976 13084
rect 4912 13024 4976 13028
rect 4992 13084 5056 13088
rect 4992 13028 4996 13084
rect 4996 13028 5052 13084
rect 5052 13028 5056 13084
rect 4992 13024 5056 13028
rect 5072 13084 5136 13088
rect 5072 13028 5076 13084
rect 5076 13028 5132 13084
rect 5132 13028 5136 13084
rect 5072 13024 5136 13028
rect 5152 13084 5216 13088
rect 5152 13028 5156 13084
rect 5156 13028 5212 13084
rect 5212 13028 5216 13084
rect 5152 13024 5216 13028
rect 5232 13084 5296 13088
rect 5232 13028 5236 13084
rect 5236 13028 5292 13084
rect 5292 13028 5296 13084
rect 5232 13024 5296 13028
rect 10912 13084 10976 13088
rect 10912 13028 10916 13084
rect 10916 13028 10972 13084
rect 10972 13028 10976 13084
rect 10912 13024 10976 13028
rect 10992 13084 11056 13088
rect 10992 13028 10996 13084
rect 10996 13028 11052 13084
rect 11052 13028 11056 13084
rect 10992 13024 11056 13028
rect 11072 13084 11136 13088
rect 11072 13028 11076 13084
rect 11076 13028 11132 13084
rect 11132 13028 11136 13084
rect 11072 13024 11136 13028
rect 11152 13084 11216 13088
rect 11152 13028 11156 13084
rect 11156 13028 11212 13084
rect 11212 13028 11216 13084
rect 11152 13024 11216 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 4912 11996 4976 12000
rect 4912 11940 4916 11996
rect 4916 11940 4972 11996
rect 4972 11940 4976 11996
rect 4912 11936 4976 11940
rect 4992 11996 5056 12000
rect 4992 11940 4996 11996
rect 4996 11940 5052 11996
rect 5052 11940 5056 11996
rect 4992 11936 5056 11940
rect 5072 11996 5136 12000
rect 5072 11940 5076 11996
rect 5076 11940 5132 11996
rect 5132 11940 5136 11996
rect 5072 11936 5136 11940
rect 5152 11996 5216 12000
rect 5152 11940 5156 11996
rect 5156 11940 5212 11996
rect 5212 11940 5216 11996
rect 5152 11936 5216 11940
rect 5232 11996 5296 12000
rect 5232 11940 5236 11996
rect 5236 11940 5292 11996
rect 5292 11940 5296 11996
rect 5232 11936 5296 11940
rect 10912 11996 10976 12000
rect 10912 11940 10916 11996
rect 10916 11940 10972 11996
rect 10972 11940 10976 11996
rect 10912 11936 10976 11940
rect 10992 11996 11056 12000
rect 10992 11940 10996 11996
rect 10996 11940 11052 11996
rect 11052 11940 11056 11996
rect 10992 11936 11056 11940
rect 11072 11996 11136 12000
rect 11072 11940 11076 11996
rect 11076 11940 11132 11996
rect 11132 11940 11136 11996
rect 11072 11936 11136 11940
rect 11152 11996 11216 12000
rect 11152 11940 11156 11996
rect 11156 11940 11212 11996
rect 11212 11940 11216 11996
rect 11152 11936 11216 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 9996 11732 10060 11796
rect 4292 11520 4356 11524
rect 4292 11464 4306 11520
rect 4306 11464 4356 11520
rect 4292 11460 4356 11464
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 4912 10908 4976 10912
rect 4912 10852 4916 10908
rect 4916 10852 4972 10908
rect 4972 10852 4976 10908
rect 4912 10848 4976 10852
rect 4992 10908 5056 10912
rect 4992 10852 4996 10908
rect 4996 10852 5052 10908
rect 5052 10852 5056 10908
rect 4992 10848 5056 10852
rect 5072 10908 5136 10912
rect 5072 10852 5076 10908
rect 5076 10852 5132 10908
rect 5132 10852 5136 10908
rect 5072 10848 5136 10852
rect 5152 10908 5216 10912
rect 5152 10852 5156 10908
rect 5156 10852 5212 10908
rect 5212 10852 5216 10908
rect 5152 10848 5216 10852
rect 5232 10908 5296 10912
rect 5232 10852 5236 10908
rect 5236 10852 5292 10908
rect 5292 10852 5296 10908
rect 5232 10848 5296 10852
rect 10912 10908 10976 10912
rect 10912 10852 10916 10908
rect 10916 10852 10972 10908
rect 10972 10852 10976 10908
rect 10912 10848 10976 10852
rect 10992 10908 11056 10912
rect 10992 10852 10996 10908
rect 10996 10852 11052 10908
rect 11052 10852 11056 10908
rect 10992 10848 11056 10852
rect 11072 10908 11136 10912
rect 11072 10852 11076 10908
rect 11076 10852 11132 10908
rect 11132 10852 11136 10908
rect 11072 10848 11136 10852
rect 11152 10908 11216 10912
rect 11152 10852 11156 10908
rect 11156 10852 11212 10908
rect 11212 10852 11216 10908
rect 11152 10848 11216 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 4912 9820 4976 9824
rect 4912 9764 4916 9820
rect 4916 9764 4972 9820
rect 4972 9764 4976 9820
rect 4912 9760 4976 9764
rect 4992 9820 5056 9824
rect 4992 9764 4996 9820
rect 4996 9764 5052 9820
rect 5052 9764 5056 9820
rect 4992 9760 5056 9764
rect 5072 9820 5136 9824
rect 5072 9764 5076 9820
rect 5076 9764 5132 9820
rect 5132 9764 5136 9820
rect 5072 9760 5136 9764
rect 5152 9820 5216 9824
rect 5152 9764 5156 9820
rect 5156 9764 5212 9820
rect 5212 9764 5216 9820
rect 5152 9760 5216 9764
rect 5232 9820 5296 9824
rect 5232 9764 5236 9820
rect 5236 9764 5292 9820
rect 5292 9764 5296 9820
rect 5232 9760 5296 9764
rect 10912 9820 10976 9824
rect 10912 9764 10916 9820
rect 10916 9764 10972 9820
rect 10972 9764 10976 9820
rect 10912 9760 10976 9764
rect 10992 9820 11056 9824
rect 10992 9764 10996 9820
rect 10996 9764 11052 9820
rect 11052 9764 11056 9820
rect 10992 9760 11056 9764
rect 11072 9820 11136 9824
rect 11072 9764 11076 9820
rect 11076 9764 11132 9820
rect 11132 9764 11136 9820
rect 11072 9760 11136 9764
rect 11152 9820 11216 9824
rect 11152 9764 11156 9820
rect 11156 9764 11212 9820
rect 11212 9764 11216 9820
rect 11152 9760 11216 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 4912 8732 4976 8736
rect 4912 8676 4916 8732
rect 4916 8676 4972 8732
rect 4972 8676 4976 8732
rect 4912 8672 4976 8676
rect 4992 8732 5056 8736
rect 4992 8676 4996 8732
rect 4996 8676 5052 8732
rect 5052 8676 5056 8732
rect 4992 8672 5056 8676
rect 5072 8732 5136 8736
rect 5072 8676 5076 8732
rect 5076 8676 5132 8732
rect 5132 8676 5136 8732
rect 5072 8672 5136 8676
rect 5152 8732 5216 8736
rect 5152 8676 5156 8732
rect 5156 8676 5212 8732
rect 5212 8676 5216 8732
rect 5152 8672 5216 8676
rect 5232 8732 5296 8736
rect 5232 8676 5236 8732
rect 5236 8676 5292 8732
rect 5292 8676 5296 8732
rect 5232 8672 5296 8676
rect 10912 8732 10976 8736
rect 10912 8676 10916 8732
rect 10916 8676 10972 8732
rect 10972 8676 10976 8732
rect 10912 8672 10976 8676
rect 10992 8732 11056 8736
rect 10992 8676 10996 8732
rect 10996 8676 11052 8732
rect 11052 8676 11056 8732
rect 10992 8672 11056 8676
rect 11072 8732 11136 8736
rect 11072 8676 11076 8732
rect 11076 8676 11132 8732
rect 11132 8676 11136 8732
rect 11072 8672 11136 8676
rect 11152 8732 11216 8736
rect 11152 8676 11156 8732
rect 11156 8676 11212 8732
rect 11212 8676 11216 8732
rect 11152 8672 11216 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 9996 7984 10060 7988
rect 9996 7928 10010 7984
rect 10010 7928 10060 7984
rect 9996 7924 10060 7928
rect 4912 7644 4976 7648
rect 4912 7588 4916 7644
rect 4916 7588 4972 7644
rect 4972 7588 4976 7644
rect 4912 7584 4976 7588
rect 4992 7644 5056 7648
rect 4992 7588 4996 7644
rect 4996 7588 5052 7644
rect 5052 7588 5056 7644
rect 4992 7584 5056 7588
rect 5072 7644 5136 7648
rect 5072 7588 5076 7644
rect 5076 7588 5132 7644
rect 5132 7588 5136 7644
rect 5072 7584 5136 7588
rect 5152 7644 5216 7648
rect 5152 7588 5156 7644
rect 5156 7588 5212 7644
rect 5212 7588 5216 7644
rect 5152 7584 5216 7588
rect 5232 7644 5296 7648
rect 5232 7588 5236 7644
rect 5236 7588 5292 7644
rect 5292 7588 5296 7644
rect 5232 7584 5296 7588
rect 10912 7644 10976 7648
rect 10912 7588 10916 7644
rect 10916 7588 10972 7644
rect 10972 7588 10976 7644
rect 10912 7584 10976 7588
rect 10992 7644 11056 7648
rect 10992 7588 10996 7644
rect 10996 7588 11052 7644
rect 11052 7588 11056 7644
rect 10992 7584 11056 7588
rect 11072 7644 11136 7648
rect 11072 7588 11076 7644
rect 11076 7588 11132 7644
rect 11132 7588 11136 7644
rect 11072 7584 11136 7588
rect 11152 7644 11216 7648
rect 11152 7588 11156 7644
rect 11156 7588 11212 7644
rect 11212 7588 11216 7644
rect 11152 7584 11216 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 4912 6556 4976 6560
rect 4912 6500 4916 6556
rect 4916 6500 4972 6556
rect 4972 6500 4976 6556
rect 4912 6496 4976 6500
rect 4992 6556 5056 6560
rect 4992 6500 4996 6556
rect 4996 6500 5052 6556
rect 5052 6500 5056 6556
rect 4992 6496 5056 6500
rect 5072 6556 5136 6560
rect 5072 6500 5076 6556
rect 5076 6500 5132 6556
rect 5132 6500 5136 6556
rect 5072 6496 5136 6500
rect 5152 6556 5216 6560
rect 5152 6500 5156 6556
rect 5156 6500 5212 6556
rect 5212 6500 5216 6556
rect 5152 6496 5216 6500
rect 5232 6556 5296 6560
rect 5232 6500 5236 6556
rect 5236 6500 5292 6556
rect 5292 6500 5296 6556
rect 5232 6496 5296 6500
rect 10912 6556 10976 6560
rect 10912 6500 10916 6556
rect 10916 6500 10972 6556
rect 10972 6500 10976 6556
rect 10912 6496 10976 6500
rect 10992 6556 11056 6560
rect 10992 6500 10996 6556
rect 10996 6500 11052 6556
rect 11052 6500 11056 6556
rect 10992 6496 11056 6500
rect 11072 6556 11136 6560
rect 11072 6500 11076 6556
rect 11076 6500 11132 6556
rect 11132 6500 11136 6556
rect 11072 6496 11136 6500
rect 11152 6556 11216 6560
rect 11152 6500 11156 6556
rect 11156 6500 11212 6556
rect 11212 6500 11216 6556
rect 11152 6496 11216 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 4912 5468 4976 5472
rect 4912 5412 4916 5468
rect 4916 5412 4972 5468
rect 4972 5412 4976 5468
rect 4912 5408 4976 5412
rect 4992 5468 5056 5472
rect 4992 5412 4996 5468
rect 4996 5412 5052 5468
rect 5052 5412 5056 5468
rect 4992 5408 5056 5412
rect 5072 5468 5136 5472
rect 5072 5412 5076 5468
rect 5076 5412 5132 5468
rect 5132 5412 5136 5468
rect 5072 5408 5136 5412
rect 5152 5468 5216 5472
rect 5152 5412 5156 5468
rect 5156 5412 5212 5468
rect 5212 5412 5216 5468
rect 5152 5408 5216 5412
rect 5232 5468 5296 5472
rect 5232 5412 5236 5468
rect 5236 5412 5292 5468
rect 5292 5412 5296 5468
rect 5232 5408 5296 5412
rect 10912 5468 10976 5472
rect 10912 5412 10916 5468
rect 10916 5412 10972 5468
rect 10972 5412 10976 5468
rect 10912 5408 10976 5412
rect 10992 5468 11056 5472
rect 10992 5412 10996 5468
rect 10996 5412 11052 5468
rect 11052 5412 11056 5468
rect 10992 5408 11056 5412
rect 11072 5468 11136 5472
rect 11072 5412 11076 5468
rect 11076 5412 11132 5468
rect 11132 5412 11136 5468
rect 11072 5408 11136 5412
rect 11152 5468 11216 5472
rect 11152 5412 11156 5468
rect 11156 5412 11212 5468
rect 11212 5412 11216 5468
rect 11152 5408 11216 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 4912 4380 4976 4384
rect 4912 4324 4916 4380
rect 4916 4324 4972 4380
rect 4972 4324 4976 4380
rect 4912 4320 4976 4324
rect 4992 4380 5056 4384
rect 4992 4324 4996 4380
rect 4996 4324 5052 4380
rect 5052 4324 5056 4380
rect 4992 4320 5056 4324
rect 5072 4380 5136 4384
rect 5072 4324 5076 4380
rect 5076 4324 5132 4380
rect 5132 4324 5136 4380
rect 5072 4320 5136 4324
rect 5152 4380 5216 4384
rect 5152 4324 5156 4380
rect 5156 4324 5212 4380
rect 5212 4324 5216 4380
rect 5152 4320 5216 4324
rect 5232 4380 5296 4384
rect 5232 4324 5236 4380
rect 5236 4324 5292 4380
rect 5292 4324 5296 4380
rect 5232 4320 5296 4324
rect 10912 4380 10976 4384
rect 10912 4324 10916 4380
rect 10916 4324 10972 4380
rect 10972 4324 10976 4380
rect 10912 4320 10976 4324
rect 10992 4380 11056 4384
rect 10992 4324 10996 4380
rect 10996 4324 11052 4380
rect 11052 4324 11056 4380
rect 10992 4320 11056 4324
rect 11072 4380 11136 4384
rect 11072 4324 11076 4380
rect 11076 4324 11132 4380
rect 11132 4324 11136 4380
rect 11072 4320 11136 4324
rect 11152 4380 11216 4384
rect 11152 4324 11156 4380
rect 11156 4324 11212 4380
rect 11212 4324 11216 4380
rect 11152 4320 11216 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 4292 3980 4356 4044
rect 10180 4040 10244 4044
rect 10180 3984 10194 4040
rect 10194 3984 10244 4040
rect 10180 3980 10244 3984
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 4912 3292 4976 3296
rect 4912 3236 4916 3292
rect 4916 3236 4972 3292
rect 4972 3236 4976 3292
rect 4912 3232 4976 3236
rect 4992 3292 5056 3296
rect 4992 3236 4996 3292
rect 4996 3236 5052 3292
rect 5052 3236 5056 3292
rect 4992 3232 5056 3236
rect 5072 3292 5136 3296
rect 5072 3236 5076 3292
rect 5076 3236 5132 3292
rect 5132 3236 5136 3292
rect 5072 3232 5136 3236
rect 5152 3292 5216 3296
rect 5152 3236 5156 3292
rect 5156 3236 5212 3292
rect 5212 3236 5216 3292
rect 5152 3232 5216 3236
rect 5232 3292 5296 3296
rect 5232 3236 5236 3292
rect 5236 3236 5292 3292
rect 5292 3236 5296 3292
rect 5232 3232 5296 3236
rect 10912 3292 10976 3296
rect 10912 3236 10916 3292
rect 10916 3236 10972 3292
rect 10972 3236 10976 3292
rect 10912 3232 10976 3236
rect 10992 3292 11056 3296
rect 10992 3236 10996 3292
rect 10996 3236 11052 3292
rect 11052 3236 11056 3292
rect 10992 3232 11056 3236
rect 11072 3292 11136 3296
rect 11072 3236 11076 3292
rect 11076 3236 11132 3292
rect 11132 3236 11136 3292
rect 11072 3232 11136 3236
rect 11152 3292 11216 3296
rect 11152 3236 11156 3292
rect 11156 3236 11212 3292
rect 11212 3236 11216 3292
rect 11152 3232 11216 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 4912 2204 4976 2208
rect 4912 2148 4916 2204
rect 4916 2148 4972 2204
rect 4972 2148 4976 2204
rect 4912 2144 4976 2148
rect 4992 2204 5056 2208
rect 4992 2148 4996 2204
rect 4996 2148 5052 2204
rect 5052 2148 5056 2204
rect 4992 2144 5056 2148
rect 5072 2204 5136 2208
rect 5072 2148 5076 2204
rect 5076 2148 5132 2204
rect 5132 2148 5136 2204
rect 5072 2144 5136 2148
rect 5152 2204 5216 2208
rect 5152 2148 5156 2204
rect 5156 2148 5212 2204
rect 5212 2148 5216 2204
rect 5152 2144 5216 2148
rect 5232 2204 5296 2208
rect 5232 2148 5236 2204
rect 5236 2148 5292 2204
rect 5292 2148 5296 2204
rect 5232 2144 5296 2148
rect 10912 2204 10976 2208
rect 10912 2148 10916 2204
rect 10916 2148 10972 2204
rect 10972 2148 10976 2204
rect 10912 2144 10976 2148
rect 10992 2204 11056 2208
rect 10992 2148 10996 2204
rect 10996 2148 11052 2204
rect 11052 2148 11056 2204
rect 10992 2144 11056 2148
rect 11072 2204 11136 2208
rect 11072 2148 11076 2204
rect 11076 2148 11132 2204
rect 11132 2148 11136 2204
rect 11072 2144 11136 2148
rect 11152 2204 11216 2208
rect 11152 2148 11156 2204
rect 11156 2148 11212 2204
rect 11212 2148 11216 2204
rect 11152 2144 11216 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
<< metal4 >>
rect 1904 14720 2304 14736
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 4904 14176 5304 14736
rect 4904 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5304 14176
rect 4904 13088 5304 14112
rect 4904 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5304 13088
rect 4904 12000 5304 13024
rect 4904 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5304 12000
rect 4291 11524 4357 11525
rect 4291 11460 4292 11524
rect 4356 11460 4357 11524
rect 4291 11459 4357 11460
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9280 2304 10304
rect 1904 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 8192 2304 9216
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 4294 4045 4354 11459
rect 4904 10912 5304 11936
rect 4904 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5304 10912
rect 4904 9824 5304 10848
rect 4904 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5304 9824
rect 4904 8736 5304 9760
rect 4904 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5304 8736
rect 4904 7648 5304 8672
rect 4904 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5304 7648
rect 4904 6560 5304 7584
rect 4904 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5304 6560
rect 4904 5472 5304 6496
rect 4904 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5304 5472
rect 4904 4384 5304 5408
rect 4904 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5304 4384
rect 4291 4044 4357 4045
rect 4291 3980 4292 4044
rect 4356 3980 4357 4044
rect 4291 3979 4357 3980
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 2752 2304 3776
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 4904 3296 5304 4320
rect 4904 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5304 3296
rect 4904 2208 5304 3232
rect 4904 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5304 2208
rect 4904 2128 5304 2144
rect 7904 14720 8304 14736
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 10904 14176 11304 14736
rect 10904 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11304 14176
rect 9995 13836 10061 13837
rect 9995 13772 9996 13836
rect 10060 13772 10061 13836
rect 9995 13771 10061 13772
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 9998 11797 10058 13771
rect 10179 13700 10245 13701
rect 10179 13636 10180 13700
rect 10244 13636 10245 13700
rect 10179 13635 10245 13636
rect 9995 11796 10061 11797
rect 9995 11732 9996 11796
rect 10060 11732 10061 11796
rect 9995 11731 10061 11732
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9280 8304 10304
rect 7904 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 8192 8304 9216
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 9998 7989 10058 11731
rect 9995 7988 10061 7989
rect 9995 7924 9996 7988
rect 10060 7924 10061 7988
rect 9995 7923 10061 7924
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 10182 4045 10242 13635
rect 10904 13088 11304 14112
rect 10904 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11304 13088
rect 10904 12000 11304 13024
rect 10904 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11304 12000
rect 10904 10912 11304 11936
rect 10904 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11304 10912
rect 10904 9824 11304 10848
rect 10904 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11304 9824
rect 10904 8736 11304 9760
rect 10904 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11304 8736
rect 10904 7648 11304 8672
rect 10904 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11304 7648
rect 10904 6560 11304 7584
rect 10904 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11304 6560
rect 10904 5472 11304 6496
rect 10904 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11304 5472
rect 10904 4384 11304 5408
rect 10904 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11304 4384
rect 10179 4044 10245 4045
rect 10179 3980 10180 4044
rect 10244 3980 10245 4044
rect 10179 3979 10245 3980
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 2752 8304 3776
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 10904 3296 11304 4320
rect 10904 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11304 3296
rect 10904 2208 11304 3232
rect 10904 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11304 2208
rect 10904 2128 11304 2144
use sky130_fd_sc_hd__buf_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_4  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _191_
timestamp 1704896540
transform -1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13064 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp 1704896540
transform -1 0 13432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9200 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9568 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_2  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _198_
timestamp 1704896540
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9384 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _200_
timestamp 1704896540
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7360 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _203_
timestamp 1704896540
transform 1 0 6992 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13708 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _207_
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _208_
timestamp 1704896540
transform -1 0 13064 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8464 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _210_
timestamp 1704896540
transform -1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5060 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1704896540
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7728 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6992 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8280 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1704896540
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1704896540
transform 1 0 6992 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _228_
timestamp 1704896540
transform 1 0 5428 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _229_
timestamp 1704896540
transform 1 0 6532 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2208 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5060 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _236_
timestamp 1704896540
transform -1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _238_
timestamp 1704896540
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _241_
timestamp 1704896540
transform 1 0 5244 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4692 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _243_
timestamp 1704896540
transform -1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _244_
timestamp 1704896540
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1704896540
transform -1 0 8096 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _246_
timestamp 1704896540
transform 1 0 6348 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6072 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _248_
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _249_
timestamp 1704896540
transform -1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10764 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _251_
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11316 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _253_
timestamp 1704896540
transform 1 0 6348 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _254_
timestamp 1704896540
transform -1 0 6992 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _255_
timestamp 1704896540
transform 1 0 6440 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _256_
timestamp 1704896540
transform -1 0 4784 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _257_
timestamp 1704896540
transform -1 0 7544 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _258_
timestamp 1704896540
transform -1 0 6808 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _260_
timestamp 1704896540
transform -1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _261_
timestamp 1704896540
transform 1 0 5796 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _262_
timestamp 1704896540
transform 1 0 6440 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _264_
timestamp 1704896540
transform -1 0 5428 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _265_
timestamp 1704896540
transform 1 0 3956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _266_
timestamp 1704896540
transform 1 0 3036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp 1704896540
transform -1 0 6256 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _268_
timestamp 1704896540
transform -1 0 5336 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _269_
timestamp 1704896540
transform 1 0 4324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _270_
timestamp 1704896540
transform -1 0 3772 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1704896540
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _272_
timestamp 1704896540
transform 1 0 3864 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _273_
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _274_
timestamp 1704896540
transform 1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _275_
timestamp 1704896540
transform 1 0 2668 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _276_
timestamp 1704896540
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1704896540
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10304 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _279_
timestamp 1704896540
transform 1 0 9016 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1704896540
transform -1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _281_
timestamp 1704896540
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _282_
timestamp 1704896540
transform 1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1704896540
transform -1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1704896540
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _286_
timestamp 1704896540
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11224 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _288_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10580 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1704896540
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1704896540
transform -1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _291_
timestamp 1704896540
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _292_
timestamp 1704896540
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _293_
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _294_
timestamp 1704896540
transform 1 0 10488 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _295_
timestamp 1704896540
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _296_
timestamp 1704896540
transform -1 0 10120 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _298_
timestamp 1704896540
transform -1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1704896540
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _301_
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _304_
timestamp 1704896540
transform -1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1704896540
transform -1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11684 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp 1704896540
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _308_
timestamp 1704896540
transform -1 0 10764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _309_
timestamp 1704896540
transform -1 0 11224 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _310_
timestamp 1704896540
transform 1 0 11224 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _312_
timestamp 1704896540
transform 1 0 12236 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _313_
timestamp 1704896540
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1704896540
transform 1 0 12328 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _316_
timestamp 1704896540
transform 1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _318_
timestamp 1704896540
transform -1 0 8096 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _319_
timestamp 1704896540
transform -1 0 7636 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _320_
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _322_
timestamp 1704896540
transform -1 0 4876 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1704896540
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _324_
timestamp 1704896540
transform -1 0 3864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _325_
timestamp 1704896540
transform 1 0 2852 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp 1704896540
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _327_
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _328_
timestamp 1704896540
transform -1 0 4324 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1704896540
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _330_
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _331_
timestamp 1704896540
transform -1 0 4232 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _332_
timestamp 1704896540
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _333_
timestamp 1704896540
transform 1 0 2852 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _334_
timestamp 1704896540
transform -1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1704896540
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _336_
timestamp 1704896540
transform 1 0 4968 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _337_
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp 1704896540
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _339_
timestamp 1704896540
transform 1 0 4968 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _340_
timestamp 1704896540
transform 1 0 5612 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp 1704896540
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _342_
timestamp 1704896540
transform 1 0 4140 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1704896540
transform -1 0 4968 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1704896540
transform -1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8096 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _346_
timestamp 1704896540
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _347_
timestamp 1704896540
transform -1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _348_
timestamp 1704896540
transform -1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _349_
timestamp 1704896540
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _350_
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _351_
timestamp 1704896540
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _352_
timestamp 1704896540
transform -1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _353_
timestamp 1704896540
transform -1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _354_
timestamp 1704896540
transform 1 0 9752 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _355_
timestamp 1704896540
transform 1 0 9660 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _356_
timestamp 1704896540
transform 1 0 8740 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _357_
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _358_
timestamp 1704896540
transform -1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _359_
timestamp 1704896540
transform 1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _360_
timestamp 1704896540
transform 1 0 11592 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _361_
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _362_
timestamp 1704896540
transform 1 0 10396 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _363_
timestamp 1704896540
transform 1 0 10672 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1704896540
transform -1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1704896540
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _367_
timestamp 1704896540
transform -1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _368_
timestamp 1704896540
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _369_
timestamp 1704896540
transform 1 0 8648 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _370_
timestamp 1704896540
transform -1 0 8924 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _371_
timestamp 1704896540
transform 1 0 1932 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _372_
timestamp 1704896540
transform 1 0 4600 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _373_
timestamp 1704896540
transform 1 0 3588 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _374_
timestamp 1704896540
transform 1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _375_
timestamp 1704896540
transform 1 0 3680 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _376_
timestamp 1704896540
transform -1 0 2576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1704896540
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1704896540
transform -1 0 4048 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1704896540
transform 1 0 7176 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1704896540
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1704896540
transform -1 0 13524 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1704896540
transform 1 0 3220 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1704896540
transform 1 0 1472 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1704896540
transform 1 0 12052 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1704896540
transform 1 0 12052 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1704896540
transform 1 0 12052 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1704896540
transform -1 0 10396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _390_
timestamp 1704896540
transform -1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1704896540
transform 1 0 12052 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1704896540
transform 1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1704896540
transform 1 0 1472 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1704896540
transform -1 0 2944 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1704896540
transform 1 0 2208 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1704896540
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1704896540
transform 1 0 2208 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1704896540
transform -1 0 6256 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1704896540
transform -1 0 7084 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1704896540
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1704896540
transform 1 0 9660 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10304 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _403_
timestamp 1704896540
transform 1 0 6440 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _404_
timestamp 1704896540
transform 1 0 4692 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1704896540
transform 1 0 12052 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1704896540
transform 1 0 7360 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1704896540
transform -1 0 10396 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1704896540
transform -1 0 2944 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1704896540
transform 1 0 1472 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1704896540
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 6440 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 6164 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 10580 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1704896540
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_67
timestamp 1704896540
transform 1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_75
timestamp 1704896540
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_106
timestamp 1704896540
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_119
timestamp 1704896540
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_127
timestamp 1704896540
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_132
timestamp 1704896540
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 1704896540
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_31
timestamp 1704896540
transform 1 0 3956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_72
timestamp 1704896540
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_76
timestamp 1704896540
transform 1 0 8096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_101
timestamp 1704896540
transform 1 0 10396 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1704896540
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_99
timestamp 1704896540
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_104
timestamp 1704896540
transform 1 0 10672 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_116
timestamp 1704896540
transform 1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_135
timestamp 1704896540
transform 1 0 13524 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_62
timestamp 1704896540
transform 1 0 6808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_74
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8556 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1704896540
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_129
timestamp 1704896540
transform 1 0 12972 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_34
timestamp 1704896540
transform 1 0 4232 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_54
timestamp 1704896540
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_66
timestamp 1704896540
transform 1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_74
timestamp 1704896540
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1704896540
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_99
timestamp 1704896540
transform 1 0 10212 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_107
timestamp 1704896540
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_112
timestamp 1704896540
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_124
timestamp 1704896540
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_136
timestamp 1704896540
transform 1 0 13616 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_30
timestamp 1704896540
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_45
timestamp 1704896540
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1704896540
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_91
timestamp 1704896540
transform 1 0 9476 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_98
timestamp 1704896540
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1704896540
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_135
timestamp 1704896540
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_36
timestamp 1704896540
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_99
timestamp 1704896540
transform 1 0 10212 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_117
timestamp 1704896540
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_135
timestamp 1704896540
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_38
timestamp 1704896540
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 1704896540
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_63
timestamp 1704896540
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_78
timestamp 1704896540
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_133
timestamp 1704896540
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_24
timestamp 1704896540
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_59
timestamp 1704896540
transform 1 0 6532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_67
timestamp 1704896540
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_99
timestamp 1704896540
transform 1 0 10212 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_123
timestamp 1704896540
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_135
timestamp 1704896540
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1704896540
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1704896540
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_65
timestamp 1704896540
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_72
timestamp 1704896540
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_83
timestamp 1704896540
transform 1 0 8740 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 1704896540
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1704896540
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_22
timestamp 1704896540
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_37
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_58
timestamp 1704896540
transform 1 0 6440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_68
timestamp 1704896540
transform 1 0 7360 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_74
timestamp 1704896540
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1704896540
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_95
timestamp 1704896540
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_99
timestamp 1704896540
transform 1 0 10212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_106
timestamp 1704896540
transform 1 0 10856 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_118
timestamp 1704896540
transform 1 0 11960 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_130
timestamp 1704896540
transform 1 0 13064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_136
timestamp 1704896540
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_90
timestamp 1704896540
transform 1 0 9384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_121
timestamp 1704896540
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_130
timestamp 1704896540
transform 1 0 13064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_136
timestamp 1704896540
transform 1 0 13616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_32
timestamp 1704896540
transform 1 0 4048 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_59
timestamp 1704896540
transform 1 0 6532 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_63
timestamp 1704896540
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_75
timestamp 1704896540
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_93
timestamp 1704896540
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_118
timestamp 1704896540
transform 1 0 11960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_135
timestamp 1704896540
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_11
timestamp 1704896540
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_18
timestamp 1704896540
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_26
timestamp 1704896540
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_38
timestamp 1704896540
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1704896540
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_68
timestamp 1704896540
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_80
timestamp 1704896540
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_102
timestamp 1704896540
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_118
timestamp 1704896540
transform 1 0 11960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_135
timestamp 1704896540
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_76
timestamp 1704896540
transform 1 0 8096 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_101
timestamp 1704896540
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_134
timestamp 1704896540
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_45
timestamp 1704896540
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_73
timestamp 1704896540
transform 1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_89
timestamp 1704896540
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_99
timestamp 1704896540
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1704896540
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_122
timestamp 1704896540
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1704896540
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_46
timestamp 1704896540
transform 1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_64
timestamp 1704896540
transform 1 0 6992 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_106
timestamp 1704896540
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_120
timestamp 1704896540
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_126
timestamp 1704896540
transform 1 0 12696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_134
timestamp 1704896540
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_62
timestamp 1704896540
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_70
timestamp 1704896540
transform 1 0 7544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_77
timestamp 1704896540
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_88
timestamp 1704896540
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_94
timestamp 1704896540
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_130
timestamp 1704896540
transform 1 0 13064 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_136
timestamp 1704896540
transform 1 0 13616 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1704896540
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_16
timestamp 1704896540
transform 1 0 2576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_24
timestamp 1704896540
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1704896540
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_43
timestamp 1704896540
transform 1 0 5060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_56
timestamp 1704896540
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_62
timestamp 1704896540
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_74
timestamp 1704896540
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1704896540
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1704896540
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_135
timestamp 1704896540
transform 1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_14
timestamp 1704896540
transform 1 0 2392 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_22
timestamp 1704896540
transform 1 0 3128 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_46
timestamp 1704896540
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1704896540
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_75
timestamp 1704896540
transform 1 0 8004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_83
timestamp 1704896540
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_90
timestamp 1704896540
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_101
timestamp 1704896540
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1704896540
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_127
timestamp 1704896540
transform 1 0 12788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_135
timestamp 1704896540
transform 1 0 13524 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_20
timestamp 1704896540
transform 1 0 2944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_117
timestamp 1704896540
transform 1 0 11868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1704896540
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_15
timestamp 1704896540
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_21
timestamp 1704896540
transform 1 0 3036 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_29
timestamp 1704896540
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1704896540
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_68
timestamp 1704896540
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_80
timestamp 1704896540
transform 1 0 8464 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_89
timestamp 1704896540
transform 1 0 9292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_101
timestamp 1704896540
transform 1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 1704896540
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_6
timestamp 1704896540
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_13
timestamp 1704896540
transform 1 0 2300 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_24
timestamp 1704896540
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_35
timestamp 1704896540
transform 1 0 4324 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_46
timestamp 1704896540
transform 1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_54
timestamp 1704896540
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_60
timestamp 1704896540
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_64
timestamp 1704896540
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_68
timestamp 1704896540
transform 1 0 7360 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 1704896540
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_90
timestamp 1704896540
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_102
timestamp 1704896540
transform 1 0 10488 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_108
timestamp 1704896540
transform 1 0 11040 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_113
timestamp 1704896540
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_119
timestamp 1704896540
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_123
timestamp 1704896540
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_135
timestamp 1704896540
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1704896540
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1704896540
transform -1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1704896540
transform -1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1704896540
transform -1 0 3680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1704896540
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1704896540
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1704896540
transform 1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1704896540
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 1704896540
transform -1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 1704896540
transform -1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1704896540
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1704896540
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 1704896540
transform -1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp 1704896540
transform -1 0 5336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1704896540
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1704896540
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output22
timestamp 1704896540
transform -1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output24
timestamp 1704896540
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 13984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 13984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 13984 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 13984 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_64
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_66
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_67
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_68
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_69
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_70
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_71
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_72
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_73
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_74
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_75
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_76
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_77
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_78
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_79
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_81
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_82
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_83
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_84
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_85
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_86
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_87
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_88
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_89
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_92
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_93
timestamp 1704896540
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_94
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_95
timestamp 1704896540
transform 1 0 11408 0 1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 4904 2128 5304 14736 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10904 2128 11304 14736 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1904 2128 2304 14736 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7904 2128 8304 14736 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 analog_comparator_out
port 2 nsew signal input
flabel metal2 s 12070 16435 12126 17235 0 FreeSans 224 90 0 0 calib_enable
port 3 nsew signal input
flabel metal2 s 14094 16435 14150 17235 0 FreeSans 224 90 0 0 clk
port 4 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 comparator_nen
port 5 nsew signal tristate
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 dac_set[0]
port 6 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 dac_set[1]
port 7 nsew signal tristate
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 dac_set[2]
port 8 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 dac_set[3]
port 9 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 dac_set[4]
port 10 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 dac_set[5]
port 11 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 dac_set[6]
port 12 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 dac_set[7]
port 13 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 do_calibrate
port 14 nsew signal tristate
flabel metal2 s 9034 16435 9090 17235 0 FreeSans 224 90 0 0 result[0]
port 15 nsew signal tristate
flabel metal2 s 8022 16435 8078 17235 0 FreeSans 224 90 0 0 result[1]
port 16 nsew signal tristate
flabel metal2 s 7010 16435 7066 17235 0 FreeSans 224 90 0 0 result[2]
port 17 nsew signal tristate
flabel metal2 s 5998 16435 6054 17235 0 FreeSans 224 90 0 0 result[3]
port 18 nsew signal tristate
flabel metal2 s 4986 16435 5042 17235 0 FreeSans 224 90 0 0 result[4]
port 19 nsew signal tristate
flabel metal2 s 3974 16435 4030 17235 0 FreeSans 224 90 0 0 result[5]
port 20 nsew signal tristate
flabel metal2 s 2962 16435 3018 17235 0 FreeSans 224 90 0 0 result[6]
port 21 nsew signal tristate
flabel metal2 s 1950 16435 2006 17235 0 FreeSans 224 90 0 0 result[7]
port 22 nsew signal tristate
flabel metal2 s 938 16435 994 17235 0 FreeSans 224 90 0 0 result_ready
port 23 nsew signal tristate
flabel metal2 s 13082 16435 13138 17235 0 FreeSans 224 90 0 0 rst
port 24 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 thresh_sel
port 25 nsew signal tristate
flabel metal2 s 10046 16435 10102 17235 0 FreeSans 224 90 0 0 use_ext_thresh
port 26 nsew signal input
flabel metal2 s 11058 16435 11114 17235 0 FreeSans 224 90 0 0 user_enable
port 27 nsew signal input
rlabel metal1 7544 14144 7544 14144 0 VGND
rlabel metal1 7544 14688 7544 14688 0 VPWR
rlabel metal1 3266 7820 3266 7820 0 _000_
rlabel metal1 3925 8534 3925 8534 0 _001_
rlabel metal1 7206 13226 7206 13226 0 _002_
rlabel metal1 6752 12818 6752 12818 0 _003_
rlabel metal1 3940 13226 3940 13226 0 _004_
rlabel metal1 3440 12818 3440 12818 0 _005_
rlabel metal2 2162 13090 2162 13090 0 _006_
rlabel metal2 12190 8738 12190 8738 0 _007_
rlabel metal1 12272 9554 12272 9554 0 _008_
rlabel metal2 10074 9826 10074 9826 0 _009_
rlabel metal1 9894 13294 9894 13294 0 _010_
rlabel viali 12369 12206 12369 12206 0 _011_
rlabel via1 10713 13226 10713 13226 0 _012_
rlabel via1 1789 5202 1789 5202 0 _013_
rlabel metal1 2806 6256 2806 6256 0 _014_
rlabel metal2 2990 5474 2990 5474 0 _015_
rlabel metal2 3726 3298 3726 3298 0 _016_
rlabel metal1 2428 3026 2428 3026 0 _017_
rlabel metal1 6036 3026 6036 3026 0 _018_
rlabel metal2 6578 3298 6578 3298 0 _019_
rlabel metal1 4692 3706 4692 3706 0 _020_
rlabel via1 9977 4114 9977 4114 0 _021_
rlabel metal1 10380 5610 10380 5610 0 _022_
rlabel metal1 6486 5066 6486 5066 0 _023_
rlabel metal1 2438 8534 2438 8534 0 _024_
rlabel via1 12369 5270 12369 5270 0 _025_
rlabel metal1 11720 4114 11720 4114 0 _026_
rlabel via1 7677 3502 7677 3502 0 _027_
rlabel metal1 9480 3026 9480 3026 0 _028_
rlabel metal2 1978 8738 1978 8738 0 _029_
rlabel metal1 1748 11322 1748 11322 0 _030_
rlabel via1 7590 8602 7590 8602 0 _031_
rlabel metal1 7498 8500 7498 8500 0 _032_
rlabel metal1 8556 5882 8556 5882 0 _033_
rlabel metal1 8694 6834 8694 6834 0 _034_
rlabel metal1 7222 8432 7222 8432 0 _035_
rlabel metal1 5796 8942 5796 8942 0 _036_
rlabel metal1 3082 13158 3082 13158 0 _037_
rlabel metal1 6486 7922 6486 7922 0 _038_
rlabel metal1 3358 9010 3358 9010 0 _039_
rlabel metal2 2990 9316 2990 9316 0 _040_
rlabel metal1 2760 9418 2760 9418 0 _041_
rlabel metal2 4002 9146 4002 9146 0 _042_
rlabel via1 5753 7854 5753 7854 0 _043_
rlabel metal2 6486 7956 6486 7956 0 _044_
rlabel metal1 6394 7514 6394 7514 0 _045_
rlabel via1 6222 7922 6222 7922 0 _046_
rlabel metal1 5014 8466 5014 8466 0 _047_
rlabel metal1 3818 8058 3818 8058 0 _048_
rlabel metal1 10442 13906 10442 13906 0 _049_
rlabel metal1 6348 9350 6348 9350 0 _050_
rlabel metal1 6486 13226 6486 13226 0 _051_
rlabel metal1 5888 11798 5888 11798 0 _052_
rlabel metal2 5106 11186 5106 11186 0 _053_
rlabel metal1 5796 11662 5796 11662 0 _054_
rlabel metal1 9568 6970 9568 6970 0 _055_
rlabel metal1 9522 11764 9522 11764 0 _056_
rlabel metal1 9154 8908 9154 8908 0 _057_
rlabel metal1 10534 7820 10534 7820 0 _058_
rlabel metal1 9246 12104 9246 12104 0 _059_
rlabel metal1 6486 13328 6486 13328 0 _060_
rlabel metal2 6854 13668 6854 13668 0 _061_
rlabel metal1 4554 11594 4554 11594 0 _062_
rlabel metal1 6762 11832 6762 11832 0 _063_
rlabel metal1 5244 12614 5244 12614 0 _064_
rlabel metal1 6026 13294 6026 13294 0 _065_
rlabel metal1 6762 13702 6762 13702 0 _066_
rlabel metal2 5750 11356 5750 11356 0 _067_
rlabel metal1 5428 10778 5428 10778 0 _068_
rlabel metal1 4278 13940 4278 13940 0 _069_
rlabel metal1 3726 13498 3726 13498 0 _070_
rlabel metal1 5520 12954 5520 12954 0 _071_
rlabel metal1 4738 13906 4738 13906 0 _072_
rlabel metal1 3358 13736 3358 13736 0 _073_
rlabel metal1 8878 9894 8878 9894 0 _074_
rlabel metal1 4508 10234 4508 10234 0 _075_
rlabel metal1 3128 11186 3128 11186 0 _076_
rlabel metal1 2254 11050 2254 11050 0 _077_
rlabel metal1 2438 11254 2438 11254 0 _078_
rlabel metal1 2392 11322 2392 11322 0 _079_
rlabel metal1 10718 9690 10718 9690 0 _080_
rlabel metal1 9660 11730 9660 11730 0 _081_
rlabel metal1 9154 9588 9154 9588 0 _082_
rlabel metal2 9706 9112 9706 9112 0 _083_
rlabel metal1 11730 8432 11730 8432 0 _084_
rlabel metal1 6578 4046 6578 4046 0 _085_
rlabel metal1 2530 8364 2530 8364 0 _086_
rlabel metal1 11960 8942 11960 8942 0 _087_
rlabel metal1 11086 9146 11086 9146 0 _088_
rlabel metal1 10166 9633 10166 9633 0 _089_
rlabel metal1 10074 9078 10074 9078 0 _090_
rlabel metal2 10810 10455 10810 10455 0 _091_
rlabel metal1 11822 10778 11822 10778 0 _092_
rlabel metal1 11040 10642 11040 10642 0 _093_
rlabel metal1 10442 10438 10442 10438 0 _094_
rlabel metal2 9614 9350 9614 9350 0 _095_
rlabel metal1 10902 12852 10902 12852 0 _096_
rlabel metal1 10212 6970 10212 6970 0 _097_
rlabel metal1 9844 12410 9844 12410 0 _098_
rlabel metal1 11546 11764 11546 11764 0 _099_
rlabel metal1 11408 12818 11408 12818 0 _100_
rlabel metal1 10396 12614 10396 12614 0 _101_
rlabel metal1 9752 12954 9752 12954 0 _102_
rlabel metal1 12558 11662 12558 11662 0 _103_
rlabel metal1 11776 11322 11776 11322 0 _104_
rlabel metal1 10994 11186 10994 11186 0 _105_
rlabel metal1 10580 11866 10580 11866 0 _106_
rlabel metal1 11546 12308 11546 12308 0 _107_
rlabel metal1 12052 11730 12052 11730 0 _108_
rlabel metal2 11224 11730 11224 11730 0 _109_
rlabel metal2 10856 13260 10856 13260 0 _110_
rlabel metal1 12604 11866 12604 11866 0 _111_
rlabel metal2 11546 13430 11546 13430 0 _112_
rlabel metal1 7222 5202 7222 5202 0 _113_
rlabel metal1 8372 5338 8372 5338 0 _114_
rlabel via1 5566 5204 5566 5204 0 _115_
rlabel metal1 5198 4488 5198 4488 0 _116_
rlabel metal1 4646 5134 4646 5134 0 _117_
rlabel metal1 2438 5644 2438 5644 0 _118_
rlabel metal1 3174 6154 3174 6154 0 _119_
rlabel metal1 3220 6290 3220 6290 0 _120_
rlabel metal1 4232 5882 4232 5882 0 _121_
rlabel metal1 3174 5236 3174 5236 0 _122_
rlabel metal1 4048 3502 4048 3502 0 _123_
rlabel metal1 3864 3026 3864 3026 0 _124_
rlabel metal2 3450 4420 3450 4420 0 _125_
rlabel metal1 1978 3604 1978 3604 0 _126_
rlabel metal1 6072 4114 6072 4114 0 _127_
rlabel metal1 7222 3502 7222 3502 0 _128_
rlabel metal1 5704 3706 5704 3706 0 _129_
rlabel metal1 6394 3094 6394 3094 0 _130_
rlabel metal2 4738 3706 4738 3706 0 _131_
rlabel metal1 4416 3502 4416 3502 0 _132_
rlabel metal1 9200 3910 9200 3910 0 _133_
rlabel metal1 10166 6834 10166 6834 0 _134_
rlabel metal1 9522 4114 9522 4114 0 _135_
rlabel metal1 9775 4590 9775 4590 0 _136_
rlabel metal1 8970 5713 8970 5713 0 _137_
rlabel metal1 9982 4624 9982 4624 0 _138_
rlabel metal1 9982 4522 9982 4522 0 _139_
rlabel metal1 8464 4590 8464 4590 0 _140_
rlabel metal1 10120 5542 10120 5542 0 _141_
rlabel metal1 7452 4590 7452 4590 0 _142_
rlabel metal1 11776 6834 11776 6834 0 _143_
rlabel metal1 10902 5032 10902 5032 0 _144_
rlabel metal1 10864 5338 10864 5338 0 _145_
rlabel metal1 11132 4590 11132 4590 0 _146_
rlabel metal1 9568 2618 9568 2618 0 _147_
rlabel metal1 8280 4114 8280 4114 0 _148_
rlabel metal1 8832 2618 8832 2618 0 _149_
rlabel metal1 8418 3060 8418 3060 0 _150_
rlabel metal2 4094 10880 4094 10880 0 _151_
rlabel metal2 3634 11220 3634 11220 0 _152_
rlabel metal2 2530 12002 2530 12002 0 _153_
rlabel metal2 3726 12104 3726 12104 0 _154_
rlabel metal1 1794 11118 1794 11118 0 _155_
rlabel metal2 9338 6698 9338 6698 0 _156_
rlabel metal1 7176 7378 7176 7378 0 _157_
rlabel metal1 6670 7174 6670 7174 0 _158_
rlabel metal1 12098 8466 12098 8466 0 _159_
rlabel metal1 11316 9554 11316 9554 0 _160_
rlabel metal1 8050 11832 8050 11832 0 _161_
rlabel metal1 6808 7922 6808 7922 0 _162_
rlabel via1 10902 12189 10902 12189 0 _163_
rlabel metal2 5934 11033 5934 11033 0 _164_
rlabel via2 6854 10659 6854 10659 0 _165_
rlabel metal1 8694 11322 8694 11322 0 _166_
rlabel metal1 7820 8058 7820 8058 0 _167_
rlabel metal1 6992 9146 6992 9146 0 _168_
rlabel metal1 6808 9622 6808 9622 0 _169_
rlabel metal1 6394 10982 6394 10982 0 _170_
rlabel metal2 12558 10574 12558 10574 0 _171_
rlabel metal1 12696 11118 12696 11118 0 _172_
rlabel metal1 4876 10642 4876 10642 0 _173_
rlabel metal1 6762 12138 6762 12138 0 _174_
rlabel metal1 8050 9996 8050 9996 0 _175_
rlabel metal1 4830 11798 4830 11798 0 _176_
rlabel metal1 6164 11594 6164 11594 0 _177_
rlabel metal1 4692 10642 4692 10642 0 _178_
rlabel metal1 4508 10778 4508 10778 0 _179_
rlabel metal2 5934 7174 5934 7174 0 _180_
rlabel metal1 10120 11730 10120 11730 0 _181_
rlabel metal1 5290 7820 5290 7820 0 _182_
rlabel metal1 11960 7378 11960 7378 0 _183_
rlabel metal1 10350 7378 10350 7378 0 _184_
rlabel metal1 10810 7786 10810 7786 0 _185_
rlabel metal2 5566 10574 5566 10574 0 _186_
rlabel metal2 7406 6086 7406 6086 0 _187_
rlabel metal2 7406 7650 7406 7650 0 _188_
rlabel metal1 13340 3706 13340 3706 0 adc.comparator.compres.ffsync.stage0
rlabel metal1 6716 6766 6716 6766 0 adc.comparator.compres.ffsync.stage1
rlabel metal1 13248 8806 13248 8806 0 adc.internalCounter\[0\]
rlabel metal1 13432 9418 13432 9418 0 adc.internalCounter\[1\]
rlabel metal1 9292 11798 9292 11798 0 adc.internalCounter\[2\]
rlabel metal1 9154 12818 9154 12818 0 adc.internalCounter\[3\]
rlabel metal1 9154 11526 9154 11526 0 adc.internalCounter\[4\]
rlabel metal1 12558 12852 12558 12852 0 adc.internalCounter\[5\]
rlabel metal1 10994 5202 10994 5202 0 adc.state\[0\]
rlabel metal1 9200 6154 9200 6154 0 adc.state\[1\]
rlabel metal1 7590 6970 7590 6970 0 adc.state\[2\]
rlabel metal1 6992 6834 6992 6834 0 adc.state\[3\]
rlabel metal1 9108 2414 9108 2414 0 adc.syncroCount\[0\]
rlabel metal1 9292 2346 9292 2346 0 adc.syncroCount\[1\]
rlabel metal2 14122 1588 14122 1588 0 analog_comparator_out
rlabel metal1 12236 14382 12236 14382 0 calib_enable
rlabel metal2 14122 12522 14122 12522 0 clk
rlabel metal1 10626 9928 10626 9928 0 clknet_0_clk
rlabel metal1 7222 3570 7222 3570 0 clknet_2_0__leaf_clk
rlabel metal1 2116 13294 2116 13294 0 clknet_2_1__leaf_clk
rlabel metal1 13432 5678 13432 5678 0 clknet_2_2__leaf_clk
rlabel metal1 12098 9588 12098 9588 0 clknet_2_3__leaf_clk
rlabel metal2 12926 959 12926 959 0 comparator_nen
rlabel metal2 966 1520 966 1520 0 dac_set[0]
rlabel metal2 2162 1520 2162 1520 0 dac_set[1]
rlabel metal2 3358 1520 3358 1520 0 dac_set[2]
rlabel metal2 4554 1520 4554 1520 0 dac_set[3]
rlabel metal2 5750 1520 5750 1520 0 dac_set[4]
rlabel metal2 6946 959 6946 959 0 dac_set[5]
rlabel metal2 8142 959 8142 959 0 dac_set[6]
rlabel metal2 9338 1656 9338 1656 0 dac_set[7]
rlabel metal2 11730 959 11730 959 0 do_calibrate
rlabel metal2 13478 3026 13478 3026 0 net1
rlabel metal1 5796 2414 5796 2414 0 net10
rlabel metal1 6187 2346 6187 2346 0 net11
rlabel metal1 8418 2448 8418 2448 0 net12
rlabel metal2 9982 2992 9982 2992 0 net13
rlabel metal1 11868 2414 11868 2414 0 net14
rlabel metal1 7640 6222 7640 6222 0 net15
rlabel metal1 7544 13974 7544 13974 0 net16
rlabel metal1 4002 5678 4002 5678 0 net17
rlabel metal1 4462 13906 4462 13906 0 net18
rlabel metal1 3312 13430 3312 13430 0 net19
rlabel metal1 12052 14246 12052 14246 0 net2
rlabel metal1 3588 7990 3588 7990 0 net20
rlabel metal2 3220 13804 3220 13804 0 net21
rlabel metal1 2530 14382 2530 14382 0 net22
rlabel metal1 1564 9146 1564 9146 0 net23
rlabel metal1 10718 2414 10718 2414 0 net24
rlabel metal1 2714 11220 2714 11220 0 net3
rlabel metal2 11408 13294 11408 13294 0 net4
rlabel metal2 13478 6052 13478 6052 0 net5
rlabel metal1 2254 2482 2254 2482 0 net6
rlabel metal1 2070 2414 2070 2414 0 net7
rlabel metal1 3726 5678 3726 5678 0 net8
rlabel metal2 4830 2587 4830 2587 0 net9
rlabel metal1 9108 14586 9108 14586 0 result[0]
rlabel metal1 8004 14586 8004 14586 0 result[1]
rlabel metal1 7084 14586 7084 14586 0 result[2]
rlabel metal1 6210 14586 6210 14586 0 result[3]
rlabel metal2 5106 15555 5106 15555 0 result[4]
rlabel metal1 4048 14586 4048 14586 0 result[5]
rlabel metal2 3082 15555 3082 15555 0 result[6]
rlabel metal1 2208 14586 2208 14586 0 result[7]
rlabel metal1 1196 14586 1196 14586 0 result_ready
rlabel metal1 13156 14382 13156 14382 0 rst
rlabel metal2 10534 959 10534 959 0 thresh_sel
rlabel metal3 10143 13668 10143 13668 0 use_ext_thresh
rlabel metal1 11132 14382 11132 14382 0 user_enable
<< properties >>
string FIXED_BBOX 0 0 15091 17235
<< end >>
