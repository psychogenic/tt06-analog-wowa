magic
tech sky130A
magscale 1 2
timestamp 1713299947
<< pwell >>
rect 5210 4190 5320 4290
rect 6200 4100 6310 4190
<< viali >>
rect 4020 6040 4070 7470
rect 3910 3790 3960 5660
rect 4820 5320 4880 7700
rect 6650 5320 6710 7700
rect 7030 4640 7070 7750
rect 4880 4220 5040 4260
rect 6510 4220 6670 4260
rect 6790 3690 6840 4010
rect 7820 3690 7870 3920
rect 8350 3690 8400 3920
rect 4010 3570 4390 3630
rect 4830 3580 6740 3630
rect 7890 3590 8330 3630
<< metal1 >>
rect 3650 7800 8500 8260
rect 3650 7790 6760 7800
rect 3650 7470 4090 7560
rect 3650 6040 4020 7470
rect 4070 6040 4090 7470
rect 4120 7010 4310 7790
rect 4550 7700 4900 7790
rect 4550 7320 4820 7700
rect 4550 7250 4610 7320
rect 4550 7190 4590 7250
rect 3650 6010 4090 6040
rect 3650 5660 3980 6010
rect 4150 5970 4520 6470
rect 3650 5620 3910 5660
rect 3650 3660 3690 5620
rect 3850 3790 3910 5620
rect 3960 3790 3980 5660
rect 4100 5520 4110 5590
rect 4290 5520 4300 5590
rect 4330 5430 4520 5970
rect 4020 5200 4520 5430
rect 4550 6330 4610 7190
rect 4550 6270 4590 6330
rect 4550 5420 4610 6270
rect 4550 5360 4590 5420
rect 4550 5330 4610 5360
rect 4780 5330 4820 7320
rect 4550 5320 4820 5330
rect 4880 5320 4900 7700
rect 5020 7650 6090 7720
rect 6290 7650 6300 7710
rect 6500 7650 6510 7710
rect 6620 7700 6760 7790
rect 5260 7640 6090 7650
rect 5260 7570 6160 7640
rect 4940 7410 6580 7570
rect 4940 7330 5660 7410
rect 5260 7320 5660 7330
rect 5030 7190 5040 7250
rect 5220 7190 5230 7250
rect 5280 7100 5660 7320
rect 4940 6850 5660 7100
rect 5260 6790 5660 6850
rect 5020 6730 5660 6790
rect 5260 6670 5660 6730
rect 4940 6430 5660 6670
rect 5030 6270 5040 6330
rect 5220 6270 5230 6330
rect 5260 6210 5660 6430
rect 4940 5970 5660 6210
rect 5260 5870 5660 5970
rect 5020 5820 5660 5870
rect 5260 5730 5660 5820
rect 4940 5490 5660 5730
rect 5030 5360 5040 5420
rect 5220 5360 5230 5420
rect 4550 5290 4900 5320
rect 5260 5280 5660 5490
rect 4330 5120 4520 5200
rect 4100 5060 4520 5120
rect 4330 4980 4520 5060
rect 4940 5040 5660 5280
rect 4020 4750 4520 4980
rect 5260 4950 5660 5040
rect 5020 4910 5660 4950
rect 5860 7330 6580 7410
rect 5860 7090 6160 7330
rect 6300 7190 6320 7250
rect 6500 7190 6510 7250
rect 5860 6850 6580 7090
rect 5860 6670 6160 6850
rect 6290 6730 6300 6790
rect 6500 6730 6510 6790
rect 5860 6430 6580 6670
rect 5860 6210 6160 6430
rect 6300 6270 6320 6330
rect 6500 6270 6510 6330
rect 5860 5970 6580 6210
rect 5860 5730 6160 5970
rect 6290 5810 6300 5870
rect 6500 5810 6510 5870
rect 5860 5490 6580 5730
rect 5860 5280 6160 5490
rect 6300 5360 6320 5420
rect 6500 5360 6510 5420
rect 6620 5320 6650 7700
rect 6710 5320 6760 7700
rect 6930 7790 8500 7800
rect 6930 7750 7080 7790
rect 6930 5870 7030 7750
rect 6940 5790 7030 5870
rect 6930 5560 7030 5790
rect 6940 5480 7030 5560
rect 6620 5290 6760 5320
rect 5860 5040 6580 5280
rect 5860 4910 6160 5040
rect 6355 4950 6465 4956
rect 5020 4900 6160 4910
rect 4100 4600 4110 4670
rect 4290 4600 4300 4670
rect 4330 4520 4520 4750
rect 5260 4720 6160 4900
rect 6290 4890 6300 4950
rect 6500 4890 6510 4950
rect 6310 4840 6355 4890
rect 6465 4840 6500 4890
rect 6355 4834 6465 4840
rect 5260 4560 5730 4720
rect 6300 4620 6310 4700
rect 4020 4290 4520 4520
rect 4680 4490 4880 4530
rect 5080 4510 5730 4560
rect 5990 4570 6310 4620
rect 6480 4570 6500 4700
rect 6710 4570 6760 5290
rect 6930 5240 7030 5480
rect 6940 4640 7030 5240
rect 7070 4640 7080 7750
rect 7210 7700 7220 7760
rect 7410 7700 7420 7760
rect 5080 4490 5540 4510
rect 5990 4500 6470 4570
rect 6710 4560 6780 4570
rect 7010 4560 7080 4640
rect 7110 5140 7180 7700
rect 7220 7540 7230 7600
rect 7420 7540 7430 7600
rect 7580 7570 8500 7610
rect 7210 7380 7220 7440
rect 7410 7380 7420 7440
rect 7220 7220 7230 7280
rect 7420 7220 7430 7280
rect 7210 7070 7220 7130
rect 7410 7070 7420 7130
rect 7220 6910 7230 6970
rect 7420 6910 7430 6970
rect 7210 6750 7220 6810
rect 7410 6750 7420 6810
rect 7220 6590 7230 6650
rect 7420 6590 7430 6650
rect 7210 6430 7220 6490
rect 7410 6430 7420 6490
rect 7220 6270 7230 6330
rect 7420 6270 7430 6330
rect 7210 6120 7220 6180
rect 7410 6120 7420 6180
rect 7220 5960 7230 6020
rect 7420 5960 7430 6020
rect 7210 5800 7220 5860
rect 7410 5800 7420 5860
rect 7220 5650 7230 5710
rect 7420 5650 7430 5710
rect 7210 5490 7220 5550
rect 7410 5490 7420 5550
rect 7220 5330 7230 5390
rect 7420 5330 7430 5390
rect 7210 5170 7220 5230
rect 7410 5170 7420 5230
rect 7110 5080 7190 5140
rect 7110 5000 7120 5080
rect 7180 5000 7190 5080
rect 7220 5010 7230 5070
rect 7420 5010 7430 5070
rect 7110 4960 7190 5000
rect 7110 4590 7180 4960
rect 7210 4850 7220 4910
rect 7410 4850 7420 4910
rect 7220 4700 7230 4760
rect 7420 4700 7430 4760
rect 7210 4540 7220 4600
rect 7410 4540 7420 4600
rect 4680 4486 4700 4490
rect 4680 4375 4695 4486
rect 4840 4452 4880 4490
rect 6650 4486 6850 4530
rect 4950 4452 4960 4470
rect 4840 4409 4960 4452
rect 4680 4370 4700 4375
rect 4840 4370 4880 4409
rect 4950 4400 4960 4409
rect 5020 4452 5030 4470
rect 5570 4452 5580 4470
rect 5020 4409 5580 4452
rect 5020 4400 5030 4409
rect 5570 4400 5580 4409
rect 5640 4400 5650 4470
rect 5870 4400 5880 4470
rect 5940 4455 5950 4470
rect 6490 4455 6500 4470
rect 5940 4410 6500 4455
rect 5940 4400 5950 4410
rect 6490 4400 6500 4410
rect 6560 4455 6570 4470
rect 6650 4455 6705 4486
rect 6560 4406 6705 4455
rect 6560 4400 6570 4406
rect 4680 4330 4880 4370
rect 6650 4376 6705 4406
rect 6815 4376 6850 4486
rect 7580 4400 7650 7570
rect 7770 7030 8390 7570
rect 8470 7030 8500 7570
rect 7770 6990 8500 7030
rect 7770 6960 8010 6990
rect 7770 4400 7840 6960
rect 8000 6930 8010 6960
rect 8200 6970 8500 6990
rect 8200 6960 8250 6970
rect 8200 6930 8210 6960
rect 8020 6920 8040 6930
rect 8030 6910 8040 6920
rect 8190 6910 8200 6930
rect 7910 6790 7980 6830
rect 7910 6600 8280 6790
rect 7910 6340 7980 6600
rect 8010 6450 8020 6510
rect 8200 6450 8210 6510
rect 8350 6500 8500 6530
rect 7910 6150 8280 6340
rect 7910 5870 7980 6150
rect 8010 5990 8020 6050
rect 8200 5990 8210 6050
rect 7910 5680 8280 5870
rect 7910 5440 7980 5680
rect 8010 5530 8020 5590
rect 8200 5530 8210 5590
rect 7910 5250 8280 5440
rect 7910 4980 7980 5250
rect 8010 5070 8020 5140
rect 8200 5070 8210 5140
rect 7910 4790 8280 4980
rect 7910 4530 7980 4790
rect 8010 4610 8020 4680
rect 8200 4610 8210 4680
rect 5090 4300 6420 4360
rect 6650 4330 6850 4376
rect 7910 4340 8280 4530
rect 5090 4290 5290 4300
rect 4330 4240 4520 4290
rect 4330 4210 4460 4240
rect 4100 4150 4460 4210
rect 4330 4110 4460 4150
rect 4590 4110 4596 4240
rect 4860 4210 4870 4270
rect 5050 4210 5060 4270
rect 5260 4160 5290 4290
rect 5370 4160 6200 4300
rect 6280 4290 6420 4300
rect 6280 4160 6310 4290
rect 6490 4210 6500 4270
rect 6680 4210 6690 4270
rect 7481 4264 7659 4270
rect 7910 4264 7980 4340
rect 4330 4070 4520 4110
rect 5260 4100 6310 4160
rect 7659 4086 7980 4264
rect 8030 4150 8040 4210
rect 8200 4150 8210 4210
rect 7481 4080 7659 4086
rect 4020 3840 4520 4070
rect 7910 4060 7980 4086
rect 3850 3660 3980 3790
rect 4330 3750 4520 3840
rect 4820 3780 4830 3960
rect 4890 3780 4900 3960
rect 4340 3740 4520 3750
rect 4990 3740 5170 4040
rect 5280 3800 5290 3940
rect 5360 3800 5370 3940
rect 5470 3740 5650 4040
rect 5740 3800 5750 3940
rect 5820 3800 5830 3940
rect 5930 3740 6110 4040
rect 6200 3800 6210 3940
rect 6280 3800 6290 3940
rect 6380 3740 6560 4040
rect 6780 4010 7050 4050
rect 6660 3780 6670 3960
rect 6730 3780 6740 3960
rect 4100 3670 4110 3740
rect 4290 3670 4300 3740
rect 4340 3680 6660 3740
rect 6780 3690 6790 4010
rect 6840 3690 7050 4010
rect 3650 3640 3980 3660
rect 6780 3640 7050 3690
rect 7540 3920 7880 3940
rect 7540 3690 7820 3920
rect 7870 3690 7880 3920
rect 7910 3870 8300 4060
rect 8350 4000 8380 6500
rect 8460 4000 8500 6500
rect 8350 3940 8500 4000
rect 8330 3920 8500 3940
rect 7910 3770 7980 3870
rect 8010 3690 8020 3760
rect 8200 3690 8210 3760
rect 8330 3690 8350 3920
rect 8400 3690 8500 3920
rect 7540 3640 7880 3690
rect 8330 3640 8500 3690
rect 3660 3630 8500 3640
rect 3660 3570 4010 3630
rect 4390 3580 4830 3630
rect 6740 3590 7890 3630
rect 8330 3590 8500 3630
rect 6740 3580 8500 3590
rect 4390 3570 8500 3580
rect 3660 3550 8500 3570
rect 3660 3400 4800 3550
rect 4900 3530 5750 3550
rect 5820 3530 6630 3550
rect 6730 3460 8500 3550
rect 6720 3400 8500 3460
rect 3660 3170 8500 3400
<< via1 >>
rect 4610 7250 4780 7320
rect 4590 7190 4780 7250
rect 3690 3660 3850 5620
rect 4110 5520 4290 5590
rect 4610 6330 4780 7190
rect 4590 6270 4780 6330
rect 4610 5420 4780 6270
rect 4590 5360 4780 5420
rect 4610 5330 4780 5360
rect 6300 7650 6500 7710
rect 5040 7190 5220 7250
rect 5040 6270 5220 6330
rect 5040 5360 5220 5420
rect 6320 7190 6500 7250
rect 6300 6730 6500 6790
rect 6320 6270 6500 6330
rect 6300 5810 6500 5870
rect 6320 5360 6500 5420
rect 6760 5870 6930 7800
rect 6760 5790 6940 5870
rect 6760 5560 6930 5790
rect 6760 5480 6940 5560
rect 4110 4600 4290 4670
rect 6300 4890 6500 4950
rect 6355 4840 6465 4890
rect 6310 4570 6480 4700
rect 6760 5240 6930 5480
rect 6760 4640 6940 5240
rect 7220 7700 7410 7760
rect 6760 4570 7010 4640
rect 6780 4560 7010 4570
rect 7230 7540 7420 7600
rect 7220 7380 7410 7440
rect 7230 7220 7420 7280
rect 7220 7070 7410 7130
rect 7230 6910 7420 6970
rect 7220 6750 7410 6810
rect 7230 6590 7420 6650
rect 7220 6430 7410 6490
rect 7230 6270 7420 6330
rect 7220 6120 7410 6180
rect 7230 5960 7420 6020
rect 7220 5800 7410 5860
rect 7230 5650 7420 5710
rect 7220 5490 7410 5550
rect 7230 5330 7420 5390
rect 7220 5170 7410 5230
rect 7120 5000 7180 5080
rect 7230 5010 7420 5070
rect 7220 4850 7410 4910
rect 7230 4700 7420 4760
rect 7220 4540 7410 4600
rect 4700 4486 4840 4490
rect 4695 4375 4840 4486
rect 4700 4370 4840 4375
rect 4960 4400 5020 4470
rect 5580 4400 5640 4470
rect 5880 4400 5940 4470
rect 6500 4400 6560 4470
rect 6705 4376 6815 4486
rect 7650 4400 7770 7570
rect 8390 7030 8470 7570
rect 8010 6930 8200 6990
rect 8040 6910 8190 6930
rect 8020 6450 8200 6510
rect 8020 5990 8200 6050
rect 8020 5530 8200 5590
rect 8020 5070 8200 5140
rect 8020 4610 8200 4680
rect 4460 4110 4590 4240
rect 4870 4260 5050 4270
rect 4870 4220 4880 4260
rect 4880 4220 5040 4260
rect 5040 4220 5050 4260
rect 4870 4210 5050 4220
rect 5290 4160 5370 4300
rect 6200 4160 6280 4300
rect 6500 4260 6680 4270
rect 6500 4220 6510 4260
rect 6510 4220 6670 4260
rect 6670 4220 6680 4260
rect 6500 4210 6680 4220
rect 7481 4086 7659 4264
rect 8040 4150 8200 4210
rect 4830 3780 4890 3960
rect 5290 3800 5360 3940
rect 5750 3800 5820 3940
rect 6210 3800 6280 3940
rect 6670 3780 6730 3960
rect 4110 3670 4290 3740
rect 8380 4000 8460 6500
rect 8020 3690 8200 3760
rect 4800 3530 4900 3550
rect 5750 3530 5820 3550
rect 6630 3530 6730 3550
rect 4800 3460 6730 3530
rect 4800 3400 6720 3460
<< metal2 >>
rect 6760 7800 6930 7810
rect 5582 7760 5938 7768
rect 5580 7710 6510 7760
rect 5582 7650 6300 7710
rect 6500 7650 6510 7710
rect 5582 7642 6500 7650
rect 4610 7320 4780 7330
rect 4590 7250 4610 7260
rect 5040 7250 5220 7260
rect 4580 7190 4590 7250
rect 4780 7190 5040 7250
rect 5220 7190 5270 7250
rect 4590 7180 4610 7190
rect 4590 6330 4610 6340
rect 5040 7180 5220 7190
rect 5582 6798 5938 7642
rect 6300 7640 6500 7642
rect 6320 7250 6760 7260
rect 6500 7190 6760 7250
rect 6320 7180 6500 7190
rect 6300 6798 6500 6800
rect 5582 6790 6510 6798
rect 5582 6730 6300 6790
rect 6500 6730 6510 6790
rect 5582 6722 6510 6730
rect 5040 6330 5220 6340
rect 4580 6270 4590 6330
rect 4780 6270 5040 6330
rect 5220 6270 5270 6330
rect 4590 6260 4610 6270
rect 3690 5620 3850 5630
rect 3850 5590 4320 5620
rect 3850 5520 4110 5590
rect 4290 5520 4320 5590
rect 3850 5490 4320 5520
rect 4590 5420 4610 5430
rect 5040 6260 5220 6270
rect 5582 5878 5938 6722
rect 6300 6720 6500 6722
rect 6320 6330 6760 6350
rect 6500 6270 6760 6330
rect 6320 6260 6500 6270
rect 6300 5878 6500 5880
rect 5582 5870 6500 5878
rect 5582 5810 6300 5870
rect 5582 5802 6500 5810
rect 5040 5420 5220 5430
rect 4580 5360 4590 5420
rect 4780 5360 5040 5420
rect 5220 5360 5270 5420
rect 4590 5350 4610 5360
rect 5040 5350 5220 5360
rect 4610 5320 4780 5330
rect 5582 5110 5938 5802
rect 6300 5800 6500 5802
rect 6930 7760 7420 7770
rect 6930 7700 7220 7760
rect 7410 7700 7420 7760
rect 6930 7690 7420 7700
rect 7220 7600 8500 7610
rect 7220 7540 7230 7600
rect 7420 7570 8500 7600
rect 7420 7540 7650 7570
rect 7220 7530 7650 7540
rect 6930 7440 7420 7450
rect 6930 7380 7220 7440
rect 7410 7380 7420 7440
rect 6930 7370 7420 7380
rect 7580 7280 7650 7530
rect 7220 7220 7230 7280
rect 7420 7220 7650 7280
rect 6930 7130 7420 7140
rect 6930 7070 7220 7130
rect 7410 7070 7420 7130
rect 6930 7060 7420 7070
rect 7580 6970 7650 7220
rect 7220 6910 7230 6970
rect 7420 6910 7650 6970
rect 6930 6810 7420 6820
rect 6930 6750 7220 6810
rect 7410 6750 7420 6810
rect 6930 6740 7420 6750
rect 7580 6650 7650 6910
rect 7220 6590 7230 6650
rect 7420 6590 7650 6650
rect 6930 6490 7410 6500
rect 6930 6430 7220 6490
rect 6930 6420 7410 6430
rect 7580 6340 7650 6590
rect 7220 6330 7650 6340
rect 7220 6270 7230 6330
rect 7420 6270 7650 6330
rect 6930 6180 7410 6190
rect 6930 6120 7220 6180
rect 6930 6110 7410 6120
rect 7580 6020 7650 6270
rect 7220 5960 7230 6020
rect 7420 5960 7650 6020
rect 7220 5950 7650 5960
rect 6940 5860 7420 5870
rect 6940 5800 7220 5860
rect 7410 5800 7420 5860
rect 6940 5790 7420 5800
rect 7580 5710 7650 5950
rect 7220 5650 7230 5710
rect 7420 5650 7650 5710
rect 7220 5640 7650 5650
rect 6940 5550 7420 5560
rect 6940 5490 7220 5550
rect 7410 5490 7420 5550
rect 6940 5480 7420 5490
rect 6320 5420 6760 5430
rect 6500 5360 6760 5420
rect 6320 5350 6500 5360
rect 5582 5102 5630 5110
rect 5584 4950 5630 5102
rect 5920 5102 5938 5110
rect 7580 5390 7650 5640
rect 7220 5330 7230 5390
rect 7420 5330 7650 5390
rect 7220 5320 7650 5330
rect 5920 4950 5936 5102
rect 6355 5065 6465 5074
rect 5584 4854 5936 4950
rect 6300 4955 6355 4960
rect 6465 4955 6500 4960
rect 6300 4950 6500 4955
rect 6300 4840 6355 4890
rect 6465 4840 6500 4890
rect 3850 4670 4320 4710
rect 3850 4600 4110 4670
rect 4290 4600 4320 4670
rect 6300 4700 6500 4840
rect 6300 4650 6310 4700
rect 3850 4580 4320 4600
rect 6480 4650 6500 4700
rect 6310 4560 6480 4570
rect 6940 5230 7420 5240
rect 6940 5170 7220 5230
rect 7410 5170 7420 5230
rect 6940 5160 7420 5170
rect 6980 5080 7180 5090
rect 7580 5080 7650 5320
rect 6980 5070 7120 5080
rect 7110 5000 7120 5070
rect 7220 5070 7650 5080
rect 7220 5010 7230 5070
rect 7420 5010 7650 5070
rect 7220 5000 7650 5010
rect 7110 4990 7180 5000
rect 6980 4980 7120 4990
rect 6940 4910 7410 4920
rect 6940 4850 7220 4910
rect 6940 4840 7410 4850
rect 7580 4770 7650 5000
rect 7220 4760 7650 4770
rect 7220 4700 7230 4760
rect 7420 4700 7650 4760
rect 7220 4690 7650 4700
rect 6940 4640 7010 4650
rect 7010 4600 7410 4620
rect 6760 4560 6780 4570
rect 7010 4560 7220 4600
rect 6990 4540 7220 4560
rect 6990 4530 7410 4540
rect 4700 4492 4840 4500
rect 4695 4490 4840 4492
rect 4695 4486 4700 4490
rect 6705 4486 6815 4492
rect 4840 4480 5635 4486
rect 5885 4480 6705 4486
rect 4840 4470 5640 4480
rect 4840 4400 4960 4470
rect 5020 4400 5580 4470
rect 4840 4390 5640 4400
rect 5880 4470 6705 4480
rect 5940 4400 6500 4470
rect 6560 4400 6705 4470
rect 5880 4390 6705 4400
rect 4840 4375 5635 4390
rect 5885 4376 6705 4390
rect 7580 4400 7650 4690
rect 7770 7030 8390 7570
rect 8470 7030 8500 7570
rect 7770 6990 8500 7030
rect 7770 6930 8010 6990
rect 8200 6970 8500 6990
rect 8200 6930 8240 6970
rect 7770 6910 8040 6930
rect 8190 6910 8240 6930
rect 7770 6880 8240 6910
rect 7770 6070 7840 6880
rect 8010 6510 8500 6530
rect 8010 6450 8020 6510
rect 8200 6500 8500 6510
rect 8200 6450 8380 6500
rect 8010 6420 8380 6450
rect 7770 6050 8240 6070
rect 7770 5990 8020 6050
rect 8200 5990 8240 6050
rect 7770 5960 8240 5990
rect 7770 5150 7840 5960
rect 8350 5620 8380 6420
rect 8010 5590 8380 5620
rect 8010 5530 8020 5590
rect 8200 5530 8380 5590
rect 8010 5510 8380 5530
rect 7770 5140 8240 5150
rect 7770 5070 8020 5140
rect 8200 5070 8240 5140
rect 7770 5040 8240 5070
rect 7770 4520 7840 5040
rect 8350 4700 8380 5510
rect 8010 4680 8380 4700
rect 8010 4610 8020 4680
rect 8200 4610 8380 4680
rect 8010 4590 8380 4610
rect 7770 4400 8200 4520
rect 4695 4370 4700 4375
rect 6705 4370 6815 4376
rect 4695 4369 4840 4370
rect 4700 4360 4840 4369
rect 5270 4300 5390 4320
rect 4790 4270 5060 4280
rect 4460 4240 4590 4246
rect 4590 4110 4595 4240
rect 4725 4110 4734 4240
rect 4790 4210 4870 4270
rect 5050 4210 5060 4270
rect 4790 4190 5060 4210
rect 4460 4104 4590 4110
rect 4790 3960 4920 4190
rect 3850 3740 4320 3790
rect 3850 3670 4110 3740
rect 4290 3670 4320 3740
rect 3850 3660 4320 3670
rect 4790 3780 4830 3960
rect 4890 3780 4920 3960
rect 3690 3650 3850 3660
rect 4790 3550 4920 3780
rect 5270 4160 5290 4300
rect 5370 4160 5390 4300
rect 5270 3940 5390 4160
rect 6180 4300 6300 4320
rect 6180 4160 6200 4300
rect 6280 4160 6300 4300
rect 7277 4290 7445 4299
rect 6480 4270 6750 4280
rect 6480 4210 6500 4270
rect 6680 4210 6750 4270
rect 6480 4190 6750 4210
rect 5270 3800 5290 3940
rect 5360 3800 5390 3940
rect 5270 3770 5390 3800
rect 5730 3940 5840 3970
rect 5730 3800 5750 3940
rect 5820 3800 5840 3940
rect 5730 3550 5840 3800
rect 6180 3940 6300 4160
rect 6180 3800 6210 3940
rect 6280 3800 6300 3940
rect 6180 3770 6300 3800
rect 6620 3960 6750 4190
rect 7272 4086 7277 4264
rect 7445 4086 7481 4264
rect 7659 4086 7665 4264
rect 8040 4210 8200 4400
rect 8040 4140 8200 4150
rect 7277 4051 7445 4060
rect 6620 3780 6670 3960
rect 6730 3780 6750 3960
rect 8350 4000 8380 4590
rect 8460 4000 8500 6500
rect 8350 3790 8500 4000
rect 6620 3550 6750 3780
rect 8010 3760 8500 3790
rect 8010 3690 8020 3760
rect 8200 3690 8500 3760
rect 8010 3680 8500 3690
rect 4790 3400 4800 3550
rect 4900 3530 5750 3550
rect 5820 3530 6630 3550
rect 6730 3460 6750 3550
rect 6720 3400 6750 3460
rect 4790 3370 6750 3400
<< via2 >>
rect 5630 4950 5920 5110
rect 6355 4955 6465 5065
rect 6980 4990 7110 5070
rect 4595 4110 4725 4240
rect 7277 4060 7445 4290
<< metal3 >>
rect 5610 5113 7000 5120
rect 5610 5110 7113 5113
rect 5610 4950 5630 5110
rect 5920 5075 7113 5110
rect 5920 5070 7120 5075
rect 5920 5065 6980 5070
rect 5920 4955 6355 5065
rect 6465 4990 6980 5065
rect 7110 4990 7120 5070
rect 6465 4985 7120 4990
rect 6465 4955 7113 4985
rect 5920 4950 7113 4955
rect 5610 4948 7113 4950
rect 5610 4930 7000 4948
rect 6070 4830 6640 4930
rect 4540 4290 7450 4295
rect 4540 4240 7277 4290
rect 4540 4110 4595 4240
rect 4725 4110 7277 4240
rect 4540 4060 7277 4110
rect 7445 4060 7450 4290
rect 4540 4055 7450 4060
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM1
timestamp 1712811291
transform 0 -1 6220 1 0 4436
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_lvt_8TELWR  XM2
timestamp 1712811291
transform 0 -1 5300 1 0 4436
box -246 -460 246 460
use sky130_fd_pr__nfet_01v8_VWWVRL  XM3
timestamp 1712811291
transform 1 0 5783 0 1 3870
box -1083 -310 1083 310
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM4
timestamp 1712811291
transform 0 1 5129 -1 0 6301
box -1541 -319 1541 319
use sky130_fd_pr__pfet_01v8_lvt_GW6ZVV  XM5
timestamp 1712811291
transform 0 -1 6399 1 0 6301
box -1541 -319 1541 319
use sky130_fd_pr__nfet_01v8_VWWVRL  XM6
timestamp 1712811291
transform 0 -1 4200 1 0 4633
box -1083 -310 1083 310
use sky130_fd_pr__nfet_01v8_WWWVRA  XM7
timestamp 1712811291
transform 0 1 8110 -1 0 5330
box -1770 -310 1770 310
use sky130_fd_pr__pfet_01v8_lvt_ER3WAW  XM8
timestamp 1712811291
transform 0 1 7319 -1 0 6147
box -1747 -319 1747 319
use sky130_fd_pr__res_xhigh_po_0p35_5BGKUX  XR1
timestamp 1712811291
transform 1 0 4201 0 1 6742
box -201 -862 201 862
<< labels >>
flabel metal1 4680 4330 4880 4530 0 FreeSans 1280 0 0 0 MINUS
port 3 nsew
flabel metal1 6650 4330 6850 4530 0 FreeSans 1280 0 0 0 PLUS
port 2 nsew
rlabel metal1 4340 5730 4510 5860 1 VBIAS
flabel metal1 7970 7240 8170 7440 0 FreeSans 1280 0 0 0 VOUT
port 4 nsew
flabel metal1 3870 3310 4070 3510 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 3980 7880 4180 8080 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
rlabel metal1 5370 4100 6200 4360 1 VX
rlabel metal3 6465 4948 6998 5113 1 V1
rlabel metal1 5260 4510 5730 4910 1 V2
rlabel space 4040 6660 4480 7400 1 V2
<< end >>
