magic
tech sky130A
magscale 1 2
timestamp 1713250549
<< pwell >>
rect 11440 7770 11520 7870
rect 16580 7650 16760 7970
rect 16730 7400 16770 7490
<< viali >>
rect 12100 10290 13700 10350
rect 14280 10220 15370 10280
rect 9790 9910 11390 9970
rect 9640 9450 9680 9840
rect 11890 9830 11940 10010
rect 11530 9560 11570 9750
rect 15980 9490 16360 9540
rect 9750 8520 9800 8910
rect 11950 8840 12000 9120
rect 13710 8580 13760 9000
rect 14130 8590 14190 9410
rect 11110 8440 11270 8480
rect 9680 7780 9720 7860
rect 10450 7580 10810 7640
rect 14170 7570 14220 7900
rect 17160 7500 17540 7550
rect 14530 7430 14910 7480
rect 16390 7430 16740 7480
rect 12760 6650 12810 6840
rect 12870 6650 12920 6840
rect 11850 6380 12660 6420
rect 13040 6380 13850 6420
<< metal1 >>
rect 9450 10720 9700 10730
rect 9450 10350 17140 10720
rect 9450 10290 12100 10350
rect 13700 10290 17140 10350
rect 9450 10280 17140 10290
rect 9450 9970 11490 10280
rect 9450 9910 9790 9970
rect 11390 9910 11490 9970
rect 9450 9900 11490 9910
rect 11675 10045 11865 10280
rect 12420 10140 12620 10230
rect 14200 10220 14280 10280
rect 15370 10220 15490 10280
rect 14200 10210 15490 10220
rect 11960 10045 12070 10050
rect 11675 10010 12070 10045
rect 9450 9840 9700 9900
rect 11675 9855 11890 10010
rect 9450 9450 9640 9840
rect 9680 9450 9700 9840
rect 11680 9830 11890 9855
rect 11940 9830 12070 10010
rect 9450 8950 9700 9450
rect 9730 9540 9820 9750
rect 9730 9220 9780 9540
rect 9820 9460 9920 9510
rect 10510 9350 10710 9830
rect 11680 9810 12070 9830
rect 14226 10114 14293 10120
rect 11680 9760 11890 9810
rect 11400 9750 11890 9760
rect 11400 9560 11530 9750
rect 11570 9560 11890 9750
rect 11400 9550 11890 9560
rect 9730 9120 9890 9220
rect 10510 9150 10760 9350
rect 10960 9150 10966 9350
rect 11680 9150 11890 9550
rect 12420 9460 12620 9940
rect 13630 10030 13740 10080
rect 14530 10110 15120 10210
rect 14226 10041 14293 10047
rect 13630 9850 13950 10030
rect 14058 9873 14283 9879
rect 13630 9840 13740 9850
rect 12781 9499 12959 9505
rect 12414 9260 12420 9460
rect 12620 9260 12626 9460
rect 12781 9315 12959 9321
rect 13771 9499 13949 9850
rect 14058 9642 14283 9648
rect 13771 9315 13949 9321
rect 14117 9640 14223 9642
rect 14117 9410 14200 9640
rect 14372 9590 14449 10060
rect 10510 9140 10710 9150
rect 11680 9120 12020 9150
rect 9450 8910 9810 8950
rect 9450 8539 9750 8910
rect 9450 8421 9451 8539
rect 9569 8520 9750 8539
rect 9800 8520 9810 8910
rect 9840 8810 9889 9120
rect 10510 9012 10710 9030
rect 9939 8849 11261 9012
rect 9840 8602 9940 8810
rect 9860 8600 9940 8602
rect 9980 8520 10074 8849
rect 10510 8830 10710 8849
rect 11098 8749 11261 8849
rect 11680 8840 11950 9120
rect 12000 8840 12020 9120
rect 11680 8815 12020 8840
rect 11690 8810 12020 8815
rect 10385 8721 10496 8727
rect 10125 8610 10385 8721
rect 10385 8604 10496 8610
rect 10780 8620 11080 8720
rect 10410 8539 10690 8550
rect 9569 8500 9810 8520
rect 9569 8421 9790 8500
rect 9450 8420 9790 8421
rect 10410 8421 10491 8539
rect 10609 8421 10690 8539
rect 9451 8415 9569 8420
rect 9460 8320 9750 8326
rect 9460 7870 9750 8118
rect 9460 7860 9840 7870
rect 9460 7780 9680 7860
rect 9720 7780 9840 7860
rect 9460 7770 9840 7780
rect 9460 6430 9750 7770
rect 10410 7690 10690 8421
rect 10780 8475 10870 8620
rect 11132 8543 11226 8749
rect 11435 8721 11546 8727
rect 11290 8620 11435 8710
rect 11546 8620 11740 8710
rect 11435 8604 11546 8610
rect 10780 8379 10870 8385
rect 11089 8480 11291 8501
rect 11425 8480 11515 8481
rect 11089 8440 11110 8480
rect 11270 8440 11291 8480
rect 11089 8320 11291 8440
rect 11420 8475 11515 8480
rect 11420 8385 11425 8475
rect 11420 8380 11515 8385
rect 11420 8340 11520 8380
rect 11089 8112 11291 8118
rect 11440 8050 11520 8340
rect 11650 8301 11740 8620
rect 11470 7870 11520 8050
rect 11440 7770 11520 7870
rect 11470 7750 11520 7770
rect 11590 8295 11760 8301
rect 11590 7780 11760 8125
rect 10410 7640 10850 7650
rect 10410 7580 10450 7640
rect 10810 7580 10850 7640
rect 10410 6430 10850 7580
rect 11590 7520 12130 7780
rect 11590 6860 11760 7520
rect 12230 7330 12450 9150
rect 12784 8760 12957 9315
rect 12510 8090 13210 8760
rect 13290 7320 13510 9140
rect 14117 9030 14130 9410
rect 13700 9000 14130 9030
rect 13700 8903 13710 9000
rect 13697 8797 13710 8903
rect 13700 8580 13710 8797
rect 13760 8590 14130 9000
rect 14190 8590 14200 9410
rect 14230 9507 14449 9590
rect 15170 9593 15247 10063
rect 15360 9990 15370 10120
rect 15450 9990 15460 10120
rect 15950 9873 16390 10280
rect 17240 10140 17440 10146
rect 17240 9934 17440 9940
rect 15792 9648 15798 9873
rect 16023 9648 16390 9873
rect 15288 9593 15294 9598
rect 15170 9510 15294 9593
rect 14230 8720 14280 9507
rect 15288 9505 15294 9510
rect 15387 9505 15393 9598
rect 15950 9540 16390 9648
rect 15950 9490 15980 9540
rect 16360 9490 16390 9540
rect 15950 9480 16390 9490
rect 16603 9609 16717 9615
rect 14470 9370 16400 9450
rect 13760 8580 14200 8590
rect 13700 8560 14200 8580
rect 14890 8510 15289 9370
rect 15410 8921 15611 8930
rect 14460 8430 15289 8510
rect 14655 8295 14825 8301
rect 14150 7900 14340 7910
rect 13580 7520 14080 7780
rect 13880 7330 14080 7520
rect 14150 7570 14170 7900
rect 14220 7650 14340 7900
rect 14220 7620 14330 7650
rect 14220 7570 14300 7620
rect 13874 7130 13880 7330
rect 14080 7130 14086 7330
rect 12220 6860 12420 7060
rect 13310 6860 13510 7050
rect 13880 6860 14080 7130
rect 11590 6660 12420 6860
rect 12220 6460 12420 6660
rect 12620 6840 13050 6860
rect 12620 6650 12760 6840
rect 12810 6650 12870 6840
rect 12920 6650 13050 6840
rect 12620 6640 13050 6650
rect 13310 6660 14080 6860
rect 12750 6430 12930 6640
rect 13310 6460 13510 6660
rect 14150 6430 14300 7570
rect 14655 7550 14825 8125
rect 15170 8020 15289 8430
rect 15409 8739 15770 8921
rect 15409 8730 15611 8739
rect 15409 8400 15591 8730
rect 15810 8510 16020 9370
rect 16603 9340 16717 9494
rect 16560 8723 16717 9340
rect 16560 8720 16650 8723
rect 15770 8430 16400 8510
rect 15410 8350 15590 8400
rect 16990 8350 17170 8356
rect 15404 8170 15410 8350
rect 15590 8170 15596 8350
rect 15130 7640 15289 8020
rect 15409 7980 15591 8170
rect 15409 7800 15780 7980
rect 15409 7799 15591 7800
rect 15151 7621 15289 7640
rect 14500 7480 14940 7500
rect 14500 7430 14530 7480
rect 14910 7430 14940 7480
rect 14500 6430 14940 7430
rect 15980 7330 16180 8120
rect 16580 7650 16770 7970
rect 16990 7880 17170 8170
rect 17250 7970 17420 9934
rect 17289 7961 17420 7970
rect 17289 7960 17867 7961
rect 17289 7910 17870 7960
rect 17289 7909 17391 7910
rect 16990 7700 17330 7880
rect 17380 7710 17640 7840
rect 17770 7710 17776 7840
rect 17810 7650 17870 7910
rect 16670 7490 16770 7650
rect 17320 7600 17870 7650
rect 15980 7124 16180 7130
rect 16330 7480 16770 7490
rect 16330 7430 16390 7480
rect 16740 7430 16770 7480
rect 16330 6430 16770 7430
rect 17130 7550 17570 7570
rect 17130 7500 17160 7550
rect 17540 7500 17570 7550
rect 17130 7476 17570 7500
rect 17130 7344 17639 7476
rect 17771 7344 17777 7476
rect 17130 6430 17570 7344
rect 9460 6420 17570 6430
rect 9460 6380 11850 6420
rect 12660 6380 13040 6420
rect 13850 6380 17570 6420
rect 9460 5990 17570 6380
<< via1 >>
rect 12420 9940 12620 10140
rect 10760 9150 10960 9350
rect 14226 10047 14293 10114
rect 12420 9260 12620 9460
rect 12781 9321 12959 9499
rect 14058 9648 14283 9873
rect 13771 9321 13949 9499
rect 9451 8421 9569 8539
rect 10385 8610 10496 8721
rect 10491 8421 10609 8539
rect 9460 8118 9750 8320
rect 11435 8610 11546 8721
rect 10780 8385 10870 8475
rect 11425 8385 11515 8475
rect 11089 8118 11291 8320
rect 11590 8125 11760 8295
rect 15370 9990 15450 10120
rect 17240 9940 17440 10140
rect 15798 9648 16023 9873
rect 15294 9505 15387 9598
rect 16603 9494 16717 9609
rect 14655 8125 14825 8295
rect 13880 7130 14080 7330
rect 15410 8170 15590 8350
rect 16990 8170 17170 8350
rect 17640 7710 17770 7840
rect 15980 7130 16180 7330
rect 17639 7344 17771 7476
<< metal2 >>
rect 12414 9940 12420 10140
rect 12620 10120 17240 10140
rect 12620 10114 15370 10120
rect 12620 10047 14226 10114
rect 14293 10047 15370 10114
rect 12620 9990 15370 10047
rect 15450 9990 17240 10120
rect 12620 9940 17240 9990
rect 17440 9940 17446 10140
rect 15798 9873 16023 9879
rect 14052 9648 14058 9873
rect 14283 9648 15798 9873
rect 15798 9642 16023 9648
rect 15283 9598 16603 9609
rect 15283 9505 15294 9598
rect 15387 9505 16603 9598
rect 12420 9460 12620 9466
rect 10760 9350 10960 9356
rect 10960 9260 12420 9350
rect 12775 9321 12781 9499
rect 12959 9321 13771 9499
rect 13949 9321 13955 9499
rect 15283 9494 16603 9505
rect 16717 9494 16723 9609
rect 10960 9150 12620 9260
rect 10760 9144 10960 9150
rect 10379 8610 10385 8721
rect 10496 8610 11435 8721
rect 11546 8610 11552 8721
rect 9445 8421 9451 8539
rect 9569 8421 10491 8539
rect 10609 8421 10615 8539
rect 10774 8385 10780 8475
rect 10870 8385 11425 8475
rect 11515 8385 11521 8475
rect 15410 8350 15590 8356
rect 9450 8320 11300 8330
rect 9450 8118 9460 8320
rect 9750 8118 11089 8320
rect 11291 8118 11300 8320
rect 11584 8125 11590 8295
rect 11760 8125 14655 8295
rect 14825 8125 14831 8295
rect 15590 8170 16990 8350
rect 17170 8170 17176 8350
rect 15410 8164 15590 8170
rect 9450 8110 11300 8118
rect 17640 7841 17770 7846
rect 17639 7840 17771 7841
rect 17639 7710 17640 7840
rect 17770 7710 17771 7840
rect 17639 7476 17771 7710
rect 17639 7338 17771 7344
rect 13880 7330 14080 7336
rect 14080 7130 15980 7330
rect 16180 7130 16186 7330
rect 13880 7124 14080 7130
use sky130_fd_pr__pfet_01v8_GGY9VD  XM1
timestamp 1712866051
transform 1 0 12856 0 1 9939
box -996 -419 996 419
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM2
timestamp 1712866051
transform 1 0 12326 0 1 8229
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM3
timestamp 1712866051
transform 1 0 13386 0 1 8229
box -396 -1019 396 1019
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM4
timestamp 1712866051
transform 1 0 13436 0 1 6760
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM5
timestamp 1712866051
transform 1 0 12246 0 1 6760
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM6
timestamp 1712866051
transform 1 0 14736 0 1 7820
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM7
timestamp 1712866051
transform 1 0 14706 0 1 8939
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM8
timestamp 1712866051
transform 1 0 16176 0 1 8939
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_UGSVTG  XM9
timestamp 1712866051
transform 0 -1 14829 1 0 10081
box -211 -719 211 719
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM10
timestamp 1712866051
transform 1 0 16176 0 1 7820
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_648S5X  XM11
timestamp 1712866051
transform 1 0 17351 0 1 7780
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_GGMWVD  XM12
timestamp 1712866051
transform 1 0 10606 0 1 9649
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM13
timestamp 1712866051
transform 1 0 10026 0 1 8709
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_lvt_FMMQLY  XM14
timestamp 1712866051
transform 1 0 11186 0 1 8670
box -296 -260 296 260
use sky130_fd_pr__nfet_01v8_lvt_FMHZDY  XM15
timestamp 1712866051
transform 1 0 10646 0 1 7820
box -996 -260 996 260
<< labels >>
rlabel metal1 15330 9380 15540 9430 1 pg2g
rlabel metal1 11590 7520 12130 7780 1 G1
rlabel metal1 9730 9120 9890 9220 1 p2p
rlabel metal2 14080 7130 15980 7330 1 G2
rlabel metal1 11440 8050 11520 8380 1 n2n
rlabel metal2 12959 9321 13771 9499 1 inhigh
rlabel metal1 14230 9507 14449 9590 1 mirhigh
flabel metal1 9850 10310 10050 10510 0 FreeSans 1280 0 0 0 VCC
port 2 nsew
flabel metal1 9800 6090 10000 6290 0 FreeSans 1280 0 0 0 VSS
port 3 nsew
flabel metal1 12240 7560 12440 7760 0 FreeSans 1280 0 0 0 MINUS
port 1 nsew
flabel metal1 13300 7560 13500 7760 0 FreeSans 1280 0 0 0 PLUS
port 0 nsew
flabel metal1 15411 8730 15611 8930 0 FreeSans 1280 0 0 0 DIFFOUT
port 6 nsew
flabel metal1 10510 8830 10710 9030 0 FreeSans 1280 0 0 0 ADJ
port 5 nsew
flabel metal1 10510 9140 10710 9340 0 FreeSans 1280 0 0 0 EN_N
port 4 nsew
<< end >>
