* NGSPICE file created from analogswitch_parax.ext - technology: sky130A

.subckt analogswitch_parax EN VCC OUT VSS IN
X0 OUT.t1 EN.t0 IN.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X1 x2.GP EN.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X2 OUT.t0 x2.GP IN.t0 VCC.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X3 VCC.t2 EN.t2 x2.GP VCC.t1 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.35
**devattr s=23200,916 d=23200,916
R0 EN EN.t0 233.88
R1 EN.n0 EN.t1 193.153
R2 EN.n0 EN.t2 174.048
R3 EN EN.n0 1.89741
R4 EN.n0 EN 1.188
R5 IN.n0 IN.t0 113.805
R6 IN IN.t1 41.5734
R7 IN.n0 IN 0.08175
R8 IN IN.n0 0.0573182
R9 OUT.n0 OUT.t0 113.803
R10 OUT OUT.t1 41.6352
R11 OUT OUT.n0 0.06925
R12 OUT.n0 OUT 0.0573182
R13 VSS.n18 VSS.n4 29056.4
R14 VSS.n9 VSS.n5 2914.44
R15 VSS.n16 VSS.n5 2914.44
R16 VSS.n16 VSS.n6 2914.44
R17 VSS.n9 VSS.n6 2914.44
R18 VSS.n21 VSS.n2 2306.06
R19 VSS.n21 VSS.n3 2306.06
R20 VSS.n23 VSS.n2 2306.06
R21 VSS.n19 VSS.n18 1994.72
R22 VSS.t0 VSS.n19 1592.68
R23 VSS.n18 VSS.n17 1159.23
R24 VSS.n22 VSS.n3 1009.07
R25 VSS.t2 VSS.n4 689.615
R26 VSS.n17 VSS.t2 689.615
R27 VSS.n3 VSS.n1 292.5
R28 VSS.n2 VSS.n0 292.5
R29 VSS.n19 VSS.n2 292.5
R30 VSS.n7 VSS.n5 292.5
R31 VSS.n5 VSS.t2 292.5
R32 VSS.n8 VSS.n6 292.5
R33 VSS.n6 VSS.t2 292.5
R34 VSS.n10 VSS.n7 189.365
R35 VSS.n15 VSS.n7 189.365
R36 VSS.n15 VSS.n14 181.929
R37 VSS.n20 VSS.n0 149.835
R38 VSS.n20 VSS.n1 149.835
R39 VSS.n24 VSS.n1 126.947
R40 VSS.n25 VSS.n0 124.462
R41 VSS.n24 VSS.n23 117.001
R42 VSS.n21 VSS.n20 117.001
R43 VSS.t0 VSS.n21 117.001
R44 VSS.n11 VSS.n10 91.8593
R45 VSS.n11 VSS.n8 85.9864
R46 VSS.n27 VSS.t1 83.7422
R47 VSS.n10 VSS.n9 73.1255
R48 VSS.n9 VSS.n4 73.1255
R49 VSS.n16 VSS.n15 73.1255
R50 VSS.n17 VSS.n16 73.1255
R51 VSS.n23 VSS.n22 62.6273
R52 VSS.n22 VSS.t0 51.1973
R53 VSS.n13 VSS.n11 9.50792
R54 VSS.n14 VSS.n13 2.3255
R55 VSS.n26 VSS.n25 1.8605
R56 VSS.n25 VSS.n24 1.2805
R57 VSS.n14 VSS.n8 0.3205
R58 VSS VSS.n12 0.315747
R59 VSS.n28 VSS 0.113
R60 VSS.n28 VSS.n27 0.0934487
R61 VSS.n26 VSS 0.088641
R62 VSS.n13 VSS 0.0518393
R63 VSS.n12 VSS 0.0402727
R64 VSS VSS.n28 0.0325513
R65 VSS.n12 VSS 0.0229359
R66 VSS.n27 VSS.n26 0.00210256
R67 VCC.n21 VCC.n15 1860
R68 VCC.n19 VCC.n18 1860
R69 VCC.n9 VCC.n3 1807.06
R70 VCC.n6 VCC.n4 1807.06
R71 VCC.n18 VCC.n17 561.481
R72 VCC.n21 VCC.n20 561.481
R73 VCC.n22 VCC.n14 198.4
R74 VCC.n16 VCC.n14 198.4
R75 VCC.n10 VCC.n2 192.754
R76 VCC.n5 VCC.n2 192.754
R77 VCC.n11 VCC.n10 183.413
R78 VCC.n9 VCC.n8 178.274
R79 VCC.n7 VCC.n6 178.274
R80 VCC.n16 VCC.n13 175.391
R81 VCC.n23 VCC.n22 173.403
R82 VCC.n25 VCC.t2 113.68
R83 VCC.n3 VCC.n1 92.5005
R84 VCC.n4 VCC.n2 92.5005
R85 VCC.n5 VCC.n0 92.2358
R86 VCC.n1 VCC.n0 87.1086
R87 VCC.n7 VCC.n3 79.3155
R88 VCC.n8 VCC.n4 79.3155
R89 VCC.n22 VCC.n21 61.6672
R90 VCC.n18 VCC.n16 61.6672
R91 VCC.n10 VCC.n9 23.1255
R92 VCC.n6 VCC.n5 23.1255
R93 VCC.n19 VCC.n14 23.1255
R94 VCC.n15 VCC.n13 23.1255
R95 VCC.n17 VCC.n15 15.947
R96 VCC.n20 VCC.n19 15.947
R97 VCC.n12 VCC.n0 9.48305
R98 VCC.t0 VCC.n7 9.12649
R99 VCC.n8 VCC.t0 9.12649
R100 VCC.n20 VCC.t1 6.98177
R101 VCC.n17 VCC.t1 6.98177
R102 VCC.n12 VCC.n11 2.3255
R103 VCC.n24 VCC.n23 1.8605
R104 VCC.n23 VCC.n13 1.0245
R105 VCC.n24 VCC 0.398648
R106 VCC.n11 VCC.n1 0.305262
R107 VCC.n26 VCC 0.124875
R108 VCC VCC.n26 0.109601
R109 VCC.n26 VCC.n25 0.105215
R110 VCC VCC.n12 0.0484167
R111 VCC.n25 VCC.n24 0.00281481
C0 EN IN 0.393415f
C1 EN x2.GP 1.13543f
C2 EN VCC 0.865357f
C3 OUT IN 0.615438f
C4 OUT x2.GP 0.235547f
C5 IN x2.GP 0.603398f
C6 OUT VCC 0.359827f
C7 IN VCC 0.302565f
C8 x2.GP VCC 1.34797f
C9 OUT EN 0.2549f
C10 EN VSS 2.52007f
C11 OUT VSS 0.789112f
C12 IN VSS 0.556176f
C13 VCC VSS 4.54035f
C14 x2.GP VSS 1.03597f
.ends

