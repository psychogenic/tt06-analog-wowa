magic
tech sky130A
magscale 1 2
timestamp 1713151418
<< metal4 >>
rect -1349 4639 1349 4680
rect -1349 2561 1093 4639
rect 1329 2561 1349 4639
rect -1349 2520 1349 2561
rect -1349 2239 1349 2280
rect -1349 161 1093 2239
rect 1329 161 1349 2239
rect -1349 120 1349 161
rect -1349 -161 1349 -120
rect -1349 -2239 1093 -161
rect 1329 -2239 1349 -161
rect -1349 -2280 1349 -2239
rect -1349 -2561 1349 -2520
rect -1349 -4639 1093 -2561
rect 1329 -4639 1349 -2561
rect -1349 -4680 1349 -4639
<< via4 >>
rect 1093 2561 1329 4639
rect 1093 161 1329 2239
rect 1093 -2239 1329 -161
rect 1093 -4639 1329 -2561
<< mimcap2 >>
rect -1269 4560 731 4600
rect -1269 2640 -1229 4560
rect 691 2640 731 4560
rect -1269 2600 731 2640
rect -1269 2160 731 2200
rect -1269 240 -1229 2160
rect 691 240 731 2160
rect -1269 200 731 240
rect -1269 -240 731 -200
rect -1269 -2160 -1229 -240
rect 691 -2160 731 -240
rect -1269 -2200 731 -2160
rect -1269 -2640 731 -2600
rect -1269 -4560 -1229 -2640
rect 691 -4560 731 -2640
rect -1269 -4600 731 -4560
<< mimcap2contact >>
rect -1229 2640 691 4560
rect -1229 240 691 2160
rect -1229 -2160 691 -240
rect -1229 -4560 691 -2640
<< metal5 >>
rect -429 4584 -109 4800
rect 1051 4639 1371 4800
rect -1253 4560 715 4584
rect -1253 2640 -1229 4560
rect 691 2640 715 4560
rect -1253 2616 715 2640
rect -429 2184 -109 2616
rect 1051 2561 1093 4639
rect 1329 2561 1371 4639
rect 1051 2239 1371 2561
rect -1253 2160 715 2184
rect -1253 240 -1229 2160
rect 691 240 715 2160
rect -1253 216 715 240
rect -429 -216 -109 216
rect 1051 161 1093 2239
rect 1329 161 1371 2239
rect 1051 -161 1371 161
rect -1253 -240 715 -216
rect -1253 -2160 -1229 -240
rect 691 -2160 715 -240
rect -1253 -2184 715 -2160
rect -429 -2616 -109 -2184
rect 1051 -2239 1093 -161
rect 1329 -2239 1371 -161
rect 1051 -2561 1371 -2239
rect -1253 -2640 715 -2616
rect -1253 -4560 -1229 -2640
rect 691 -4560 715 -2640
rect -1253 -4584 715 -4560
rect -429 -4800 -109 -4584
rect 1051 -4639 1093 -2561
rect 1329 -4639 1371 -2561
rect 1051 -4800 1371 -4639
<< properties >>
string FIXED_BBOX -1349 2520 811 4680
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
