magic
tech sky130A
magscale 1 2
timestamp 1713490400
<< viali >>
rect 1409 14569 1443 14603
rect 2145 14569 2179 14603
rect 3157 14569 3191 14603
rect 4169 14569 4203 14603
rect 5181 14569 5215 14603
rect 6377 14569 6411 14603
rect 7205 14569 7239 14603
rect 8217 14569 8251 14603
rect 9229 14569 9263 14603
rect 1593 14365 1627 14399
rect 2329 14365 2363 14399
rect 3341 14365 3375 14399
rect 4353 14365 4387 14399
rect 5365 14365 5399 14399
rect 6561 14365 6595 14399
rect 7389 14365 7423 14399
rect 8401 14365 8435 14399
rect 9413 14365 9447 14399
rect 11713 14365 11747 14399
rect 12449 14365 12483 14399
rect 13461 14365 13495 14399
rect 11529 14229 11563 14263
rect 12265 14229 12299 14263
rect 13369 14229 13403 14263
rect 3157 13889 3191 13923
rect 4261 13889 4295 13923
rect 6653 13889 6687 13923
rect 6745 13889 6779 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 7297 13889 7331 13923
rect 9689 13889 9723 13923
rect 9873 13889 9907 13923
rect 10241 13889 10275 13923
rect 3249 13821 3283 13855
rect 3709 13821 3743 13855
rect 3433 13753 3467 13787
rect 2973 13685 3007 13719
rect 4077 13685 4111 13719
rect 6377 13685 6411 13719
rect 7205 13685 7239 13719
rect 10149 13685 10183 13719
rect 3433 13481 3467 13515
rect 5457 13481 5491 13515
rect 8493 13481 8527 13515
rect 5365 13413 5399 13447
rect 2053 13277 2087 13311
rect 3985 13277 4019 13311
rect 4252 13277 4286 13311
rect 6837 13277 6871 13311
rect 7113 13277 7147 13311
rect 9413 13277 9447 13311
rect 11538 13277 11572 13311
rect 11805 13277 11839 13311
rect 11897 13277 11931 13311
rect 2320 13209 2354 13243
rect 6570 13209 6604 13243
rect 7380 13209 7414 13243
rect 12164 13209 12198 13243
rect 9229 13141 9263 13175
rect 10425 13141 10459 13175
rect 13277 13141 13311 13175
rect 2237 12937 2271 12971
rect 4445 12937 4479 12971
rect 5365 12937 5399 12971
rect 6929 12937 6963 12971
rect 7665 12937 7699 12971
rect 8953 12937 8987 12971
rect 11161 12937 11195 12971
rect 10517 12869 10551 12903
rect 12265 12869 12299 12903
rect 2053 12801 2087 12835
rect 2329 12801 2363 12835
rect 2596 12801 2630 12835
rect 4629 12801 4663 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 6653 12801 6687 12835
rect 6745 12801 6779 12835
rect 7021 12801 7055 12835
rect 7205 12801 7239 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 8033 12801 8067 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 8677 12801 8711 12835
rect 8861 12801 8895 12835
rect 10066 12801 10100 12835
rect 10425 12801 10459 12835
rect 10701 12801 10735 12835
rect 10977 12801 11011 12835
rect 11253 12801 11287 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12081 12801 12115 12835
rect 4169 12733 4203 12767
rect 4261 12733 4295 12767
rect 4537 12733 4571 12767
rect 4813 12733 4847 12767
rect 4905 12733 4939 12767
rect 4997 12733 5031 12767
rect 5089 12733 5123 12767
rect 5825 12733 5859 12767
rect 8401 12733 8435 12767
rect 8493 12733 8527 12767
rect 10333 12733 10367 12767
rect 11805 12733 11839 12767
rect 11897 12733 11931 12767
rect 5273 12665 5307 12699
rect 5457 12665 5491 12699
rect 7849 12665 7883 12699
rect 3709 12597 3743 12631
rect 3985 12597 4019 12631
rect 10885 12597 10919 12631
rect 10977 12597 11011 12631
rect 2513 12393 2547 12427
rect 3801 12393 3835 12427
rect 4537 12393 4571 12427
rect 5457 12393 5491 12427
rect 6469 12393 6503 12427
rect 7389 12393 7423 12427
rect 7849 12393 7883 12427
rect 10241 12393 10275 12427
rect 12081 12393 12115 12427
rect 2697 12325 2731 12359
rect 3065 12325 3099 12359
rect 8125 12325 8159 12359
rect 11069 12325 11103 12359
rect 11897 12325 11931 12359
rect 12817 12325 12851 12359
rect 3525 12257 3559 12291
rect 4997 12257 5031 12291
rect 3249 12189 3283 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4445 12189 4479 12223
rect 4721 12189 4755 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5733 12189 5767 12223
rect 5825 12189 5859 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 6653 12189 6687 12223
rect 7481 12189 7515 12223
rect 7757 12189 7791 12223
rect 8217 12189 8251 12223
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 9493 12189 9527 12223
rect 9689 12189 9723 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 10057 12189 10091 12223
rect 10609 12189 10643 12223
rect 10701 12189 10735 12223
rect 10793 12189 10827 12223
rect 11253 12189 11287 12223
rect 11529 12189 11563 12223
rect 11713 12189 11747 12223
rect 11805 12189 11839 12223
rect 12173 12189 12207 12223
rect 12265 12189 12299 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 12725 12199 12759 12233
rect 12909 12189 12943 12223
rect 2973 12121 3007 12155
rect 4353 12121 4387 12155
rect 6837 12121 6871 12155
rect 10977 12121 11011 12155
rect 11437 12121 11471 12155
rect 12357 12121 12391 12155
rect 4169 12053 4203 12087
rect 9413 12053 9447 12087
rect 10425 12053 10459 12087
rect 12455 12053 12489 12087
rect 3065 11849 3099 11883
rect 3525 11849 3559 11883
rect 4537 11849 4571 11883
rect 7113 11849 7147 11883
rect 7849 11849 7883 11883
rect 9965 11849 9999 11883
rect 10241 11849 10275 11883
rect 12081 11849 12115 11883
rect 3341 11713 3375 11747
rect 4721 11713 4755 11747
rect 4997 11713 5031 11747
rect 5181 11713 5215 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 7757 11713 7791 11747
rect 7849 11713 7883 11747
rect 9689 11713 9723 11747
rect 10057 11713 10091 11747
rect 10241 11713 10275 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 12440 11713 12474 11747
rect 3249 11645 3283 11679
rect 3617 11645 3651 11679
rect 3709 11645 3743 11679
rect 7481 11645 7515 11679
rect 8125 11645 8159 11679
rect 9965 11645 9999 11679
rect 11621 11645 11655 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 7941 11577 7975 11611
rect 9781 11509 9815 11543
rect 13553 11509 13587 11543
rect 1501 11305 1535 11339
rect 7389 11305 7423 11339
rect 10149 11305 10183 11339
rect 11345 11305 11379 11339
rect 12817 11305 12851 11339
rect 13185 11305 13219 11339
rect 2881 11169 2915 11203
rect 10885 11169 10919 11203
rect 11437 11169 11471 11203
rect 3157 11101 3191 11135
rect 3433 11101 3467 11135
rect 3617 11101 3651 11135
rect 4353 11101 4387 11135
rect 4813 11101 4847 11135
rect 4997 11101 5031 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 7205 11101 7239 11135
rect 7389 11101 7423 11135
rect 10057 11101 10091 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 10425 11101 10459 11135
rect 10977 11101 11011 11135
rect 11069 11101 11103 11135
rect 11161 11101 11195 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 12817 11101 12851 11135
rect 12909 11101 12943 11135
rect 2636 11033 2670 11067
rect 2973 11033 3007 11067
rect 4721 11033 4755 11067
rect 12449 11033 12483 11067
rect 4905 10965 4939 10999
rect 6561 10965 6595 10999
rect 9781 10965 9815 10999
rect 10333 10965 10367 10999
rect 12725 10965 12759 10999
rect 3525 10761 3559 10795
rect 4721 10761 4755 10795
rect 7573 10761 7607 10795
rect 7665 10761 7699 10795
rect 8493 10761 8527 10795
rect 9781 10761 9815 10795
rect 9873 10761 9907 10795
rect 10517 10761 10551 10795
rect 11069 10761 11103 10795
rect 12265 10761 12299 10795
rect 12633 10761 12667 10795
rect 12817 10693 12851 10727
rect 3157 10625 3191 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 4905 10625 4939 10659
rect 5181 10625 5215 10659
rect 5365 10625 5399 10659
rect 5825 10625 5859 10659
rect 6469 10625 6503 10659
rect 6929 10625 6963 10659
rect 7389 10625 7423 10659
rect 7757 10625 7791 10659
rect 7941 10625 7975 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 9689 10625 9723 10659
rect 10149 10625 10183 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 11713 10625 11747 10659
rect 12357 10625 12391 10659
rect 12725 10625 12759 10659
rect 2973 10557 3007 10591
rect 3065 10557 3099 10591
rect 3249 10557 3283 10591
rect 3433 10557 3467 10591
rect 3893 10557 3927 10591
rect 5917 10557 5951 10591
rect 6561 10557 6595 10591
rect 6745 10557 6779 10591
rect 8125 10557 8159 10591
rect 10241 10557 10275 10591
rect 11989 10557 12023 10591
rect 12449 10557 12483 10591
rect 12633 10557 12667 10591
rect 3801 10489 3835 10523
rect 4997 10489 5031 10523
rect 5089 10489 5123 10523
rect 6193 10489 6227 10523
rect 9505 10489 9539 10523
rect 10057 10489 10091 10523
rect 5825 10421 5859 10455
rect 7113 10421 7147 10455
rect 10149 10421 10183 10455
rect 11805 10421 11839 10455
rect 4813 10217 4847 10251
rect 9413 10217 9447 10251
rect 12173 10217 12207 10251
rect 3433 10081 3467 10115
rect 6929 10081 6963 10115
rect 7573 10081 7607 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 8585 10081 8619 10115
rect 10333 10081 10367 10115
rect 3157 10013 3191 10047
rect 3249 10013 3283 10047
rect 3341 10013 3375 10047
rect 4261 10013 4295 10047
rect 6653 10013 6687 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 7711 10013 7745 10047
rect 8033 10013 8067 10047
rect 8401 10013 8435 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9505 10013 9539 10047
rect 9781 10013 9815 10047
rect 9873 10013 9907 10047
rect 10057 10013 10091 10047
rect 4445 9945 4479 9979
rect 6285 9945 6319 9979
rect 10425 9945 10459 9979
rect 10701 9945 10735 9979
rect 2973 9877 3007 9911
rect 4077 9877 4111 9911
rect 6469 9877 6503 9911
rect 6745 9877 6779 9911
rect 7297 9877 7331 9911
rect 7849 9877 7883 9911
rect 9045 9877 9079 9911
rect 9229 9877 9263 9911
rect 3249 9673 3283 9707
rect 4169 9673 4203 9707
rect 4629 9673 4663 9707
rect 8493 9673 8527 9707
rect 9045 9673 9079 9707
rect 11529 9605 11563 9639
rect 11713 9605 11747 9639
rect 11897 9605 11931 9639
rect 2053 9537 2087 9571
rect 3433 9537 3467 9571
rect 4353 9537 4387 9571
rect 4629 9537 4663 9571
rect 4997 9537 5031 9571
rect 5365 9537 5399 9571
rect 5825 9537 5859 9571
rect 5917 9537 5951 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 7205 9537 7239 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7573 9537 7607 9571
rect 8254 9537 8288 9571
rect 8401 9537 8435 9571
rect 8861 9537 8895 9571
rect 8953 9537 8987 9571
rect 9137 9537 9171 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 10978 9527 11012 9561
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 2145 9469 2179 9503
rect 2605 9469 2639 9503
rect 2789 9469 2823 9503
rect 2973 9469 3007 9503
rect 3065 9469 3099 9503
rect 3341 9469 3375 9503
rect 3801 9469 3835 9503
rect 3985 9469 4019 9503
rect 4077 9469 4111 9503
rect 4445 9469 4479 9503
rect 8033 9469 8067 9503
rect 8769 9469 8803 9503
rect 2329 9401 2363 9435
rect 5549 9401 5583 9435
rect 9873 9401 9907 9435
rect 11253 9401 11287 9435
rect 1869 9333 1903 9367
rect 6929 9333 6963 9367
rect 7757 9333 7791 9367
rect 8125 9333 8159 9367
rect 8677 9333 8711 9367
rect 11989 9333 12023 9367
rect 2881 9129 2915 9163
rect 5365 9129 5399 9163
rect 6377 9129 6411 9163
rect 7573 9129 7607 9163
rect 7941 9129 7975 9163
rect 9045 9129 9079 9163
rect 10425 9129 10459 9163
rect 10977 9129 11011 9163
rect 11897 9129 11931 9163
rect 3893 9061 3927 9095
rect 5273 9061 5307 9095
rect 9321 9061 9355 9095
rect 11253 9061 11287 9095
rect 3157 8993 3191 9027
rect 3617 8993 3651 9027
rect 4077 8993 4111 9027
rect 12173 8993 12207 9027
rect 1501 8925 1535 8959
rect 3249 8925 3283 8959
rect 4169 8925 4203 8959
rect 4537 8925 4571 8959
rect 4629 8925 4663 8959
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 5017 8925 5051 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6561 8925 6595 8959
rect 6837 8925 6871 8959
rect 6938 8925 6972 8959
rect 7297 8925 7331 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9505 8925 9539 8959
rect 10550 8925 10584 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 11621 8925 11655 8959
rect 11713 8925 11747 8959
rect 12429 8925 12463 8959
rect 1768 8857 1802 8891
rect 6193 8857 6227 8891
rect 7113 8857 7147 8891
rect 7481 8857 7515 8891
rect 11989 8857 12023 8891
rect 2973 8789 3007 8823
rect 3433 8789 3467 8823
rect 3525 8789 3559 8823
rect 4353 8789 4387 8823
rect 4445 8789 4479 8823
rect 5825 8789 5859 8823
rect 10609 8789 10643 8823
rect 13553 8789 13587 8823
rect 4261 8585 4295 8619
rect 4445 8585 4479 8619
rect 8033 8585 8067 8619
rect 3249 8517 3283 8551
rect 9321 8517 9355 8551
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 7205 8449 7239 8483
rect 10425 8449 10459 8483
rect 12817 8449 12851 8483
rect 3341 8381 3375 8415
rect 3893 8381 3927 8415
rect 4077 8381 4111 8415
rect 4169 8381 4203 8415
rect 4905 8381 4939 8415
rect 4997 8381 5031 8415
rect 5089 8381 5123 8415
rect 2973 8313 3007 8347
rect 3617 8313 3651 8347
rect 10517 8313 10551 8347
rect 2789 8245 2823 8279
rect 3801 8245 3835 8279
rect 4629 8245 4663 8279
rect 7021 8245 7055 8279
rect 12633 8245 12667 8279
rect 7757 8041 7791 8075
rect 8125 8041 8159 8075
rect 8953 8041 8987 8075
rect 10517 8041 10551 8075
rect 11529 8041 11563 8075
rect 12265 8041 12299 8075
rect 12449 8041 12483 8075
rect 11253 7973 11287 8007
rect 8493 7905 8527 7939
rect 12173 7905 12207 7939
rect 12633 7905 12667 7939
rect 2789 7837 2823 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 11713 7837 11747 7871
rect 11897 7837 11931 7871
rect 12449 7837 12483 7871
rect 9137 7769 9171 7803
rect 9321 7769 9355 7803
rect 10701 7769 10735 7803
rect 11253 7769 11287 7803
rect 12909 7769 12943 7803
rect 2605 7701 2639 7735
rect 4353 7701 4387 7735
rect 8401 7701 8435 7735
rect 10333 7701 10367 7735
rect 10793 7701 10827 7735
rect 11805 7701 11839 7735
rect 9045 7497 9079 7531
rect 10425 7497 10459 7531
rect 13461 7497 13495 7531
rect 2320 7429 2354 7463
rect 3709 7361 3743 7395
rect 7021 7361 7055 7395
rect 8217 7361 8251 7395
rect 8401 7361 8435 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9505 7361 9539 7395
rect 10149 7361 10183 7395
rect 11069 7361 11103 7395
rect 11529 7361 11563 7395
rect 12081 7361 12115 7395
rect 12541 7361 12575 7395
rect 12909 7361 12943 7395
rect 13277 7361 13311 7395
rect 2053 7293 2087 7327
rect 7297 7293 7331 7327
rect 8493 7293 8527 7327
rect 10425 7293 10459 7327
rect 11345 7293 11379 7327
rect 3433 7225 3467 7259
rect 8217 7225 8251 7259
rect 11805 7225 11839 7259
rect 3525 7157 3559 7191
rect 6837 7157 6871 7191
rect 7205 7157 7239 7191
rect 9321 7157 9355 7191
rect 10241 7157 10275 7191
rect 5457 6953 5491 6987
rect 8125 6953 8159 6987
rect 9321 6953 9355 6987
rect 9505 6953 9539 6987
rect 10425 6953 10459 6987
rect 10517 6953 10551 6987
rect 13093 6953 13127 6987
rect 9873 6885 9907 6919
rect 10793 6885 10827 6919
rect 4077 6817 4111 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 4344 6749 4378 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 6193 6749 6227 6783
rect 8033 6749 8067 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 9137 6749 9171 6783
rect 9510 6749 9544 6783
rect 9689 6749 9723 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11345 6749 11379 6783
rect 11444 6749 11478 6783
rect 12909 6749 12943 6783
rect 6009 6681 6043 6715
rect 6438 6681 6472 6715
rect 8953 6681 8987 6715
rect 11704 6681 11738 6715
rect 7573 6613 7607 6647
rect 12817 6613 12851 6647
rect 4169 6409 4203 6443
rect 11897 6409 11931 6443
rect 3056 6341 3090 6375
rect 6009 6341 6043 6375
rect 7389 6341 7423 6375
rect 8125 6341 8159 6375
rect 8309 6341 8343 6375
rect 2329 6273 2363 6307
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 7200 6273 7234 6307
rect 7297 6273 7331 6307
rect 7572 6273 7606 6307
rect 7665 6273 7699 6307
rect 8401 6273 8435 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8769 6273 8803 6307
rect 8953 6273 8987 6307
rect 9413 6273 9447 6307
rect 9597 6273 9631 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 10701 6273 10735 6307
rect 11161 6273 11195 6307
rect 12081 6273 12115 6307
rect 12541 6273 12575 6307
rect 2789 6205 2823 6239
rect 10793 6205 10827 6239
rect 12265 6205 12299 6239
rect 6653 6137 6687 6171
rect 7941 6137 7975 6171
rect 11069 6137 11103 6171
rect 2053 6069 2087 6103
rect 4721 6069 4755 6103
rect 7021 6069 7055 6103
rect 9137 6069 9171 6103
rect 9229 6069 9263 6103
rect 9505 6069 9539 6103
rect 10425 6069 10459 6103
rect 10885 6069 10919 6103
rect 11253 6069 11287 6103
rect 12081 6069 12115 6103
rect 3065 5865 3099 5899
rect 9137 5865 9171 5899
rect 10057 5797 10091 5831
rect 10149 5797 10183 5831
rect 5457 5729 5491 5763
rect 9229 5729 9263 5763
rect 1593 5661 1627 5695
rect 1860 5661 1894 5695
rect 3249 5661 3283 5695
rect 3525 5661 3559 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 7113 5661 7147 5695
rect 7297 5661 7331 5695
rect 9505 5661 9539 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 10517 5661 10551 5695
rect 5365 5593 5399 5627
rect 5702 5593 5736 5627
rect 2973 5525 3007 5559
rect 3433 5525 3467 5559
rect 3801 5525 3835 5559
rect 4169 5525 4203 5559
rect 6837 5525 6871 5559
rect 6929 5525 6963 5559
rect 8953 5525 8987 5559
rect 9781 5525 9815 5559
rect 11805 5525 11839 5559
rect 9774 5321 9808 5355
rect 10425 5321 10459 5355
rect 12909 5321 12943 5355
rect 2636 5253 2670 5287
rect 2973 5253 3007 5287
rect 11774 5253 11808 5287
rect 2881 5185 2915 5219
rect 3249 5185 3283 5219
rect 3341 5185 3375 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 4353 5185 4387 5219
rect 4445 5185 4479 5219
rect 4629 5185 4663 5219
rect 6653 5185 6687 5219
rect 9321 5185 9355 5219
rect 9505 5185 9539 5219
rect 9597 5185 9631 5219
rect 9689 5185 9723 5219
rect 9873 5185 9907 5219
rect 9965 5185 9999 5219
rect 10609 5185 10643 5219
rect 10793 5185 10827 5219
rect 10241 5117 10275 5151
rect 10701 5117 10735 5151
rect 10885 5117 10919 5151
rect 11529 5117 11563 5151
rect 10057 5049 10091 5083
rect 10149 5049 10183 5083
rect 1501 4981 1535 5015
rect 3985 4981 4019 5015
rect 6469 4981 6503 5015
rect 9505 4981 9539 5015
rect 9321 4777 9355 4811
rect 9689 4777 9723 4811
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 4445 4573 4479 4607
rect 5089 4573 5123 4607
rect 5181 4573 5215 4607
rect 5273 4573 5307 4607
rect 5457 4573 5491 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 9873 4573 9907 4607
rect 10057 4573 10091 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 10425 4573 10459 4607
rect 13553 4573 13587 4607
rect 13308 4505 13342 4539
rect 4721 4437 4755 4471
rect 4813 4437 4847 4471
rect 10609 4437 10643 4471
rect 12173 4437 12207 4471
rect 6377 4233 6411 4267
rect 13553 4233 13587 4267
rect 3792 4165 3826 4199
rect 7573 4165 7607 4199
rect 8217 4165 8251 4199
rect 3065 4097 3099 4131
rect 3157 4097 3191 4131
rect 3249 4097 3283 4131
rect 3433 4097 3467 4131
rect 5457 4097 5491 4131
rect 5641 4097 5675 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 6561 4097 6595 4131
rect 6745 4097 6779 4131
rect 6837 4097 6871 4131
rect 7849 4097 7883 4131
rect 8033 4097 8067 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 8861 4097 8895 4131
rect 9137 4097 9171 4131
rect 9321 4097 9355 4131
rect 10221 4097 10255 4131
rect 12173 4097 12207 4131
rect 12440 4097 12474 4131
rect 3525 4029 3559 4063
rect 8585 4029 8619 4063
rect 9965 4029 9999 4063
rect 7941 3961 7975 3995
rect 9321 3961 9355 3995
rect 2789 3893 2823 3927
rect 4905 3893 4939 3927
rect 6101 3893 6135 3927
rect 7481 3893 7515 3927
rect 7757 3893 7791 3927
rect 9045 3893 9079 3927
rect 11345 3893 11379 3927
rect 4353 3689 4387 3723
rect 5825 3689 5859 3723
rect 11805 3689 11839 3723
rect 4445 3553 4479 3587
rect 2237 3485 2271 3519
rect 3893 3485 3927 3519
rect 4169 3485 4203 3519
rect 5917 3485 5951 3519
rect 6184 3485 6218 3519
rect 7389 3485 7423 3519
rect 8953 3485 8987 3519
rect 10425 3485 10459 3519
rect 10692 3485 10726 3519
rect 2504 3417 2538 3451
rect 3985 3417 4019 3451
rect 4712 3417 4746 3451
rect 7656 3417 7690 3451
rect 9198 3417 9232 3451
rect 3617 3349 3651 3383
rect 7297 3349 7331 3383
rect 8769 3349 8803 3383
rect 10333 3349 10367 3383
rect 3065 3145 3099 3179
rect 3433 3145 3467 3179
rect 6377 3145 6411 3179
rect 6745 3145 6779 3179
rect 8677 3145 8711 3179
rect 8953 3145 8987 3179
rect 4874 3077 4908 3111
rect 8493 3077 8527 3111
rect 3249 3009 3283 3043
rect 3525 3009 3559 3043
rect 4629 3009 4663 3043
rect 6561 3009 6595 3043
rect 6834 3031 6868 3065
rect 8769 3009 8803 3043
rect 8861 3009 8895 3043
rect 9965 3009 9999 3043
rect 10241 3009 10275 3043
rect 8493 2873 8527 2907
rect 6009 2805 6043 2839
rect 10425 2805 10459 2839
rect 4997 2601 5031 2635
rect 13553 2601 13587 2635
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 3985 2397 4019 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 5365 2397 5399 2431
rect 5457 2397 5491 2431
rect 6101 2397 6135 2431
rect 7297 2397 7331 2431
rect 8493 2397 8527 2431
rect 9689 2397 9723 2431
rect 10885 2397 10919 2431
rect 12081 2397 12115 2431
rect 13277 2397 13311 2431
rect 13737 2397 13771 2431
rect 1409 2261 1443 2295
rect 2329 2261 2363 2295
rect 3801 2261 3835 2295
rect 4721 2261 4755 2295
rect 5917 2261 5951 2295
rect 7113 2261 7147 2295
rect 8309 2261 8343 2295
rect 9505 2261 9539 2295
rect 10701 2261 10735 2295
rect 11897 2261 11931 2295
rect 13093 2261 13127 2295
<< metal1 >>
rect 1104 14714 14076 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 14076 14714
rect 1104 14640 14076 14662
rect 1026 14560 1032 14612
rect 1084 14600 1090 14612
rect 1397 14603 1455 14609
rect 1397 14600 1409 14603
rect 1084 14572 1409 14600
rect 1084 14560 1090 14572
rect 1397 14569 1409 14572
rect 1443 14569 1455 14603
rect 1397 14563 1455 14569
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2314 14600 2320 14612
rect 2179 14572 2320 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 3108 14572 3157 14600
rect 3108 14560 3114 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 4120 14572 4169 14600
rect 4120 14560 4126 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 5132 14572 5181 14600
rect 5132 14560 5138 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 6086 14560 6092 14612
rect 6144 14600 6150 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 6144 14572 6377 14600
rect 6144 14560 6150 14572
rect 6365 14569 6377 14572
rect 6411 14569 6423 14603
rect 6365 14563 6423 14569
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 7156 14572 7205 14600
rect 7156 14560 7162 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7892 14572 8217 14600
rect 7892 14560 7898 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 9180 14572 9229 14600
rect 9180 14560 9186 14572
rect 9217 14569 9229 14572
rect 9263 14569 9275 14603
rect 9217 14563 9275 14569
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 2498 14396 2504 14408
rect 2363 14368 2504 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 1596 14328 1624 14359
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 3510 14396 3516 14408
rect 3375 14368 3516 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 4338 14356 4344 14408
rect 4396 14356 4402 14408
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 5353 14399 5411 14405
rect 5353 14396 5365 14399
rect 4488 14368 5365 14396
rect 4488 14356 4494 14368
rect 5353 14365 5365 14368
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 5776 14368 6561 14396
rect 5776 14356 5782 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7377 14399 7435 14405
rect 7377 14396 7389 14399
rect 6972 14368 7389 14396
rect 6972 14356 6978 14368
rect 7377 14365 7389 14368
rect 7423 14365 7435 14399
rect 7377 14359 7435 14365
rect 8386 14356 8392 14408
rect 8444 14356 8450 14408
rect 9398 14356 9404 14408
rect 9456 14356 9462 14408
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 11204 14368 11713 14396
rect 11204 14356 11210 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12216 14368 12449 14396
rect 12216 14356 12222 14368
rect 12437 14365 12449 14368
rect 12483 14365 12495 14399
rect 12437 14359 12495 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 13228 14368 13461 14396
rect 13228 14356 13234 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 5442 14328 5448 14340
rect 1596 14300 5448 14328
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 12250 14220 12256 14272
rect 12308 14220 12314 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13357 14263 13415 14269
rect 13357 14260 13369 14263
rect 13320 14232 13369 14260
rect 13320 14220 13326 14232
rect 13357 14229 13369 14232
rect 13403 14229 13415 14263
rect 13357 14223 13415 14229
rect 1104 14170 14076 14192
rect 1104 14118 4918 14170
rect 4970 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 5238 14170
rect 5290 14118 10918 14170
rect 10970 14118 10982 14170
rect 11034 14118 11046 14170
rect 11098 14118 11110 14170
rect 11162 14118 11174 14170
rect 11226 14118 11238 14170
rect 11290 14118 14076 14170
rect 1104 14096 14076 14118
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13920 4307 13923
rect 5350 13920 5356 13932
rect 4295 13892 5356 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 3160 13852 3188 13883
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 5500 13892 6653 13920
rect 5500 13880 5506 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 6822 13880 6828 13932
rect 6880 13880 6886 13932
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 9674 13880 9680 13932
rect 9732 13880 9738 13932
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9824 13892 9873 13920
rect 9824 13880 9830 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10275 13892 10732 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 3160 13824 3249 13852
rect 3237 13821 3249 13824
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 10704 13796 10732 13892
rect 3421 13787 3479 13793
rect 3421 13753 3433 13787
rect 3467 13784 3479 13787
rect 4522 13784 4528 13796
rect 3467 13756 4528 13784
rect 3467 13753 3479 13756
rect 3421 13747 3479 13753
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 5316 13756 9444 13784
rect 5316 13744 5322 13756
rect 9416 13728 9444 13756
rect 10686 13744 10692 13796
rect 10744 13744 10750 13796
rect 2958 13676 2964 13728
rect 3016 13676 3022 13728
rect 4065 13719 4123 13725
rect 4065 13685 4077 13719
rect 4111 13716 4123 13719
rect 4154 13716 4160 13728
rect 4111 13688 4160 13716
rect 4111 13685 4123 13688
rect 4065 13679 4123 13685
rect 4154 13676 4160 13688
rect 4212 13676 4218 13728
rect 6362 13676 6368 13728
rect 6420 13676 6426 13728
rect 7190 13676 7196 13728
rect 7248 13676 7254 13728
rect 9398 13676 9404 13728
rect 9456 13676 9462 13728
rect 10137 13719 10195 13725
rect 10137 13685 10149 13719
rect 10183 13716 10195 13719
rect 11330 13716 11336 13728
rect 10183 13688 11336 13716
rect 10183 13685 10195 13688
rect 10137 13679 10195 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 1104 13626 14076 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 14076 13626
rect 1104 13552 14076 13574
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 5258 13512 5264 13524
rect 3476 13484 5264 13512
rect 3476 13472 3482 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5442 13472 5448 13524
rect 5500 13472 5506 13524
rect 8386 13512 8392 13524
rect 5920 13484 8392 13512
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 5353 13447 5411 13453
rect 5353 13444 5365 13447
rect 5040 13416 5365 13444
rect 5040 13404 5046 13416
rect 5353 13413 5365 13416
rect 5399 13444 5411 13447
rect 5920 13444 5948 13484
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 9674 13512 9680 13524
rect 8536 13484 9680 13512
rect 8536 13472 8542 13484
rect 9674 13472 9680 13484
rect 9732 13512 9738 13524
rect 9950 13512 9956 13524
rect 9732 13484 9956 13512
rect 9732 13472 9738 13484
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 5399 13416 5948 13444
rect 5399 13413 5411 13416
rect 5353 13407 5411 13413
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2130 13308 2136 13320
rect 2087 13280 2136 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 2866 13308 2872 13320
rect 2188 13280 2872 13308
rect 2188 13268 2194 13280
rect 2866 13268 2872 13280
rect 2924 13308 2930 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 2924 13280 3985 13308
rect 2924 13268 2930 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4240 13311 4298 13317
rect 4240 13277 4252 13311
rect 4286 13277 4298 13311
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 4240 13271 4298 13277
rect 4356 13280 6837 13308
rect 2314 13249 2320 13252
rect 2308 13203 2320 13249
rect 2314 13200 2320 13203
rect 2372 13200 2378 13252
rect 3988 13172 4016 13271
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4264 13240 4292 13271
rect 4212 13212 4292 13240
rect 4212 13200 4218 13212
rect 4356 13172 4384 13280
rect 6825 13277 6837 13280
rect 6871 13308 6883 13311
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6871 13280 7113 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 9401 13311 9459 13317
rect 9401 13277 9413 13311
rect 9447 13308 9459 13311
rect 9674 13308 9680 13320
rect 9447 13280 9680 13308
rect 9447 13277 9459 13280
rect 9401 13271 9459 13277
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 11526 13311 11584 13317
rect 11526 13308 11538 13311
rect 10376 13280 11538 13308
rect 10376 13268 10382 13280
rect 11526 13277 11538 13280
rect 11572 13277 11584 13311
rect 11526 13271 11584 13277
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11839 13280 11897 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 11885 13277 11897 13280
rect 11931 13308 11943 13311
rect 11931 13280 12296 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12268 13252 12296 13280
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 6558 13243 6616 13249
rect 6558 13240 6570 13243
rect 6420 13212 6570 13240
rect 6420 13200 6426 13212
rect 6558 13209 6570 13212
rect 6604 13209 6616 13243
rect 6558 13203 6616 13209
rect 7368 13243 7426 13249
rect 7368 13209 7380 13243
rect 7414 13240 7426 13243
rect 7650 13240 7656 13252
rect 7414 13212 7656 13240
rect 7414 13209 7426 13212
rect 7368 13203 7426 13209
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 10226 13240 10232 13252
rect 8352 13212 10232 13240
rect 8352 13200 8358 13212
rect 10226 13200 10232 13212
rect 10284 13240 10290 13252
rect 12152 13243 12210 13249
rect 10284 13212 10824 13240
rect 10284 13200 10290 13212
rect 3988 13144 4384 13172
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 6914 13172 6920 13184
rect 5500 13144 6920 13172
rect 5500 13132 5506 13144
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 9214 13132 9220 13184
rect 9272 13132 9278 13184
rect 10413 13175 10471 13181
rect 10413 13141 10425 13175
rect 10459 13172 10471 13175
rect 10686 13172 10692 13184
rect 10459 13144 10692 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10796 13172 10824 13212
rect 12152 13209 12164 13243
rect 12198 13209 12210 13243
rect 12152 13203 12210 13209
rect 11606 13172 11612 13184
rect 10796 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12176 13172 12204 13203
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 12124 13144 12204 13172
rect 12124 13132 12130 13144
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 13265 13175 13323 13181
rect 13265 13172 13277 13175
rect 12400 13144 13277 13172
rect 12400 13132 12406 13144
rect 13265 13141 13277 13144
rect 13311 13141 13323 13175
rect 13265 13135 13323 13141
rect 1104 13082 14076 13104
rect 1104 13030 4918 13082
rect 4970 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 5238 13082
rect 5290 13030 10918 13082
rect 10970 13030 10982 13082
rect 11034 13030 11046 13082
rect 11098 13030 11110 13082
rect 11162 13030 11174 13082
rect 11226 13030 11238 13082
rect 11290 13030 14076 13082
rect 1104 13008 14076 13030
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2314 12968 2320 12980
rect 2271 12940 2320 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4479 12940 4936 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4908 12912 4936 12940
rect 5350 12928 5356 12980
rect 5408 12928 5414 12980
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7098 12968 7104 12980
rect 6963 12940 7104 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 7650 12928 7656 12980
rect 7708 12928 7714 12980
rect 8941 12971 8999 12977
rect 8941 12937 8953 12971
rect 8987 12968 8999 12971
rect 9674 12968 9680 12980
rect 8987 12940 9680 12968
rect 8987 12937 8999 12940
rect 8941 12931 8999 12937
rect 9674 12928 9680 12940
rect 9732 12968 9738 12980
rect 11149 12971 11207 12977
rect 11149 12968 11161 12971
rect 9732 12940 10548 12968
rect 9732 12928 9738 12940
rect 2130 12860 2136 12912
rect 2188 12900 2194 12912
rect 2188 12872 2360 12900
rect 2188 12860 2194 12872
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12832 2099 12835
rect 2222 12832 2228 12844
rect 2087 12804 2228 12832
rect 2087 12801 2099 12804
rect 2041 12795 2099 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2332 12841 2360 12872
rect 4890 12860 4896 12912
rect 4948 12860 4954 12912
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2584 12835 2642 12841
rect 2584 12801 2596 12835
rect 2630 12832 2642 12835
rect 2958 12832 2964 12844
rect 2630 12804 2964 12832
rect 2630 12801 2642 12804
rect 2584 12795 2642 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 4617 12835 4675 12841
rect 4080 12804 4292 12832
rect 4080 12776 4108 12804
rect 4062 12724 4068 12776
rect 4120 12724 4126 12776
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 4264 12773 4292 12804
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 6365 12835 6423 12841
rect 4663 12804 5120 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 4571 12736 4660 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 4632 12708 4660 12736
rect 4798 12724 4804 12776
rect 4856 12724 4862 12776
rect 4890 12724 4896 12776
rect 4948 12724 4954 12776
rect 5092 12773 5120 12804
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12733 5043 12767
rect 4985 12727 5043 12733
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5166 12764 5172 12776
rect 5123 12736 5172 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 5000 12696 5028 12727
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 5813 12727 5871 12733
rect 4672 12668 5028 12696
rect 5261 12699 5319 12705
rect 4672 12656 4678 12668
rect 5261 12665 5273 12699
rect 5307 12696 5319 12699
rect 5445 12699 5503 12705
rect 5445 12696 5457 12699
rect 5307 12668 5457 12696
rect 5307 12665 5319 12668
rect 5261 12659 5319 12665
rect 5445 12665 5457 12668
rect 5491 12665 5503 12699
rect 5445 12659 5503 12665
rect 3326 12588 3332 12640
rect 3384 12628 3390 12640
rect 3697 12631 3755 12637
rect 3697 12628 3709 12631
rect 3384 12600 3709 12628
rect 3384 12588 3390 12600
rect 3697 12597 3709 12600
rect 3743 12628 3755 12631
rect 3786 12628 3792 12640
rect 3743 12600 3792 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 5828 12628 5856 12727
rect 4019 12600 5856 12628
rect 6380 12628 6408 12795
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 6914 12832 6920 12844
rect 6779 12804 6920 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 6656 12764 6684 12795
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7208 12841 7236 12928
rect 9214 12900 9220 12912
rect 7300 12872 8524 12900
rect 7300 12844 7328 12872
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 8021 12835 8079 12841
rect 7423 12804 7880 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7392 12764 7420 12795
rect 6656 12736 7420 12764
rect 7024 12708 7052 12736
rect 7006 12656 7012 12708
rect 7064 12656 7070 12708
rect 7852 12705 7880 12804
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12665 7895 12699
rect 7837 12659 7895 12665
rect 6822 12628 6828 12640
rect 6380 12600 6828 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 6822 12588 6828 12600
rect 6880 12628 6886 12640
rect 7650 12628 7656 12640
rect 6880 12600 7656 12628
rect 6880 12588 6886 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8036 12628 8064 12795
rect 8128 12696 8156 12795
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 8386 12724 8392 12776
rect 8444 12724 8450 12776
rect 8496 12773 8524 12872
rect 8680 12872 9220 12900
rect 8680 12841 8708 12872
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 9858 12900 9864 12912
rect 9364 12872 9864 12900
rect 9364 12860 9370 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 10520 12909 10548 12940
rect 10796 12940 11161 12968
rect 10505 12903 10563 12909
rect 10008 12872 10456 12900
rect 10008 12860 10014 12872
rect 10428 12841 10456 12872
rect 10505 12869 10517 12903
rect 10551 12900 10563 12903
rect 10551 12872 10640 12900
rect 10551 12869 10563 12872
rect 10505 12863 10563 12869
rect 10612 12844 10640 12872
rect 10796 12844 10824 12940
rect 11149 12937 11161 12940
rect 11195 12937 11207 12971
rect 11149 12931 11207 12937
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11296 12940 11836 12968
rect 11296 12928 11302 12940
rect 11330 12900 11336 12912
rect 11256 12872 11336 12900
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12832 8907 12835
rect 10054 12835 10112 12841
rect 10054 12832 10066 12835
rect 8895 12804 10066 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 10054 12801 10066 12804
rect 10100 12801 10112 12835
rect 10054 12795 10112 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10594 12792 10600 12844
rect 10652 12792 10658 12844
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 11256 12841 11284 12872
rect 11330 12860 11336 12872
rect 11388 12860 11394 12912
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12801 11299 12835
rect 11241 12795 11299 12801
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 9306 12764 9312 12776
rect 8527 12736 9312 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 9122 12696 9128 12708
rect 8128 12668 9128 12696
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 10336 12696 10364 12727
rect 10502 12724 10508 12776
rect 10560 12764 10566 12776
rect 10980 12764 11008 12795
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 11701 12835 11759 12841
rect 11701 12834 11713 12835
rect 11624 12806 11713 12834
rect 11624 12776 11652 12806
rect 11701 12801 11713 12806
rect 11747 12801 11759 12835
rect 11808 12832 11836 12940
rect 12066 12928 12072 12980
rect 12124 12928 12130 12980
rect 12084 12900 12112 12928
rect 12253 12903 12311 12909
rect 12253 12900 12265 12903
rect 12084 12872 12265 12900
rect 12253 12869 12265 12872
rect 12299 12869 12311 12903
rect 12253 12863 12311 12869
rect 12066 12832 12072 12844
rect 11808 12804 12072 12832
rect 11701 12795 11759 12801
rect 12066 12792 12072 12804
rect 12124 12832 12130 12844
rect 12342 12832 12348 12844
rect 12124 12804 12348 12832
rect 12124 12792 12130 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 10560 12736 11008 12764
rect 10560 12724 10566 12736
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 11882 12724 11888 12776
rect 11940 12764 11946 12776
rect 12710 12764 12716 12776
rect 11940 12736 12716 12764
rect 11940 12724 11946 12736
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 12158 12696 12164 12708
rect 10336 12668 12164 12696
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 8478 12628 8484 12640
rect 8036 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10778 12628 10784 12640
rect 9732 12600 10784 12628
rect 9732 12588 9738 12600
rect 10778 12588 10784 12600
rect 10836 12628 10842 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10836 12600 10885 12628
rect 10836 12588 10842 12600
rect 10873 12597 10885 12600
rect 10919 12597 10931 12631
rect 10873 12591 10931 12597
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12628 11023 12631
rect 11238 12628 11244 12640
rect 11011 12600 11244 12628
rect 11011 12597 11023 12600
rect 10965 12591 11023 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 12250 12628 12256 12640
rect 11388 12600 12256 12628
rect 11388 12588 11394 12600
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 12526 12628 12532 12640
rect 12308 12600 12532 12628
rect 12308 12588 12314 12600
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 1104 12538 14076 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 14076 12538
rect 1104 12464 14076 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2501 12427 2559 12433
rect 2501 12424 2513 12427
rect 2372 12396 2513 12424
rect 2372 12384 2378 12396
rect 2501 12393 2513 12396
rect 2547 12393 2559 12427
rect 2501 12387 2559 12393
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3752 12396 3801 12424
rect 3752 12384 3758 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 4522 12384 4528 12436
rect 4580 12384 4586 12436
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5224 12396 5457 12424
rect 5224 12384 5230 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5445 12387 5503 12393
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 6546 12424 6552 12436
rect 6503 12396 6552 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 2685 12359 2743 12365
rect 2685 12325 2697 12359
rect 2731 12356 2743 12359
rect 3053 12359 3111 12365
rect 3053 12356 3065 12359
rect 2731 12328 3065 12356
rect 2731 12325 2743 12328
rect 2685 12319 2743 12325
rect 3053 12325 3065 12328
rect 3099 12325 3111 12359
rect 3053 12319 3111 12325
rect 3418 12316 3424 12368
rect 3476 12316 3482 12368
rect 4890 12356 4896 12368
rect 3620 12328 4896 12356
rect 3436 12288 3464 12316
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 3160 12260 3372 12288
rect 3436 12260 3525 12288
rect 2958 12112 2964 12164
rect 3016 12112 3022 12164
rect 3160 12084 3188 12260
rect 3344 12229 3372 12260
rect 3513 12257 3525 12260
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3620 12232 3648 12328
rect 4890 12316 4896 12328
rect 4948 12356 4954 12368
rect 5350 12356 5356 12368
rect 4948 12328 5356 12356
rect 4948 12316 4954 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5552 12328 5948 12356
rect 5552 12300 5580 12328
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 3844 12260 4997 12288
rect 3844 12248 3850 12260
rect 4985 12257 4997 12260
rect 5031 12288 5043 12291
rect 5442 12288 5448 12300
rect 5031 12260 5448 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5534 12248 5540 12300
rect 5592 12248 5598 12300
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3602 12220 3608 12232
rect 3467 12192 3608 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3252 12152 3280 12183
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 3878 12180 3884 12232
rect 3936 12180 3942 12232
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4246 12180 4252 12232
rect 4304 12180 4310 12232
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4522 12220 4528 12232
rect 4479 12192 4528 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4522 12180 4528 12192
rect 4580 12220 4586 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4580 12192 4721 12220
rect 4580 12180 4586 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 3896 12152 3924 12180
rect 3252 12124 3924 12152
rect 3988 12152 4016 12180
rect 4264 12152 4292 12180
rect 3988 12124 4292 12152
rect 4341 12155 4399 12161
rect 4341 12121 4353 12155
rect 4387 12152 4399 12155
rect 4816 12152 4844 12183
rect 4890 12180 4896 12232
rect 4948 12180 4954 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5534 12152 5540 12164
rect 4387 12124 5540 12152
rect 4387 12121 4399 12124
rect 4341 12115 4399 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 5736 12152 5764 12183
rect 5810 12180 5816 12232
rect 5868 12180 5874 12232
rect 5920 12229 5948 12328
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6472 12220 6500 12387
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 6788 12396 7389 12424
rect 6788 12384 6794 12396
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 8386 12424 8392 12436
rect 7883 12396 8392 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10318 12424 10324 12436
rect 10275 12396 10324 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10410 12384 10416 12436
rect 10468 12424 10474 12436
rect 10468 12396 11100 12424
rect 10468 12384 10474 12396
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 8113 12359 8171 12365
rect 8113 12356 8125 12359
rect 6972 12328 8125 12356
rect 6972 12316 6978 12328
rect 8113 12325 8125 12328
rect 8159 12325 8171 12359
rect 8113 12319 8171 12325
rect 10778 12316 10784 12368
rect 10836 12316 10842 12368
rect 11072 12365 11100 12396
rect 11606 12384 11612 12436
rect 11664 12384 11670 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 11756 12396 12081 12424
rect 11756 12384 11762 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 12069 12387 12127 12393
rect 12167 12396 12940 12424
rect 11057 12359 11115 12365
rect 11057 12325 11069 12359
rect 11103 12325 11115 12359
rect 11057 12319 11115 12325
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11514 12356 11520 12368
rect 11296 12328 11520 12356
rect 11296 12316 11302 12328
rect 10134 12288 10140 12300
rect 7484 12260 10140 12288
rect 6135 12192 6500 12220
rect 6641 12223 6699 12229
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7006 12220 7012 12232
rect 6687 12192 7012 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6656 12152 6684 12183
rect 7006 12180 7012 12192
rect 7064 12220 7070 12232
rect 7484 12229 7512 12260
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10796 12288 10824 12316
rect 11348 12288 11376 12328
rect 11514 12316 11520 12328
rect 11572 12316 11578 12368
rect 11624 12356 11652 12384
rect 11624 12328 11836 12356
rect 11808 12288 11836 12328
rect 11882 12316 11888 12368
rect 11940 12316 11946 12368
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 12167 12356 12195 12396
rect 12805 12359 12863 12365
rect 12805 12356 12817 12359
rect 12032 12328 12195 12356
rect 12268 12328 12817 12356
rect 12032 12316 12038 12328
rect 12268 12288 12296 12328
rect 12805 12325 12817 12328
rect 12851 12325 12863 12359
rect 12805 12319 12863 12325
rect 10796 12260 11284 12288
rect 11348 12260 11652 12288
rect 11808 12260 12296 12288
rect 7469 12223 7527 12229
rect 7064 12192 7328 12220
rect 7064 12180 7070 12192
rect 7300 12164 7328 12192
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7616 12192 7757 12220
rect 7616 12180 7622 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 7745 12183 7803 12189
rect 8128 12192 8217 12220
rect 5736 12124 6684 12152
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12121 6883 12155
rect 6825 12115 6883 12121
rect 3694 12084 3700 12096
rect 3160 12056 3700 12084
rect 3694 12044 3700 12056
rect 3752 12084 3758 12096
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 3752 12056 4169 12084
rect 3752 12044 3758 12056
rect 4157 12053 4169 12056
rect 4203 12084 4215 12087
rect 4614 12084 4620 12096
rect 4203 12056 4620 12084
rect 4203 12053 4215 12056
rect 4157 12047 4215 12053
rect 4614 12044 4620 12056
rect 4672 12084 4678 12096
rect 4890 12084 4896 12096
rect 4672 12056 4896 12084
rect 4672 12044 4678 12056
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 6840 12084 6868 12115
rect 7282 12112 7288 12164
rect 7340 12112 7346 12164
rect 8128 12096 8156 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8478 12180 8484 12232
rect 8536 12220 8542 12232
rect 9033 12223 9091 12229
rect 9033 12220 9045 12223
rect 8536 12192 9045 12220
rect 8536 12180 8542 12192
rect 9033 12189 9045 12192
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9481 12223 9539 12229
rect 9481 12220 9493 12223
rect 9324 12192 9493 12220
rect 9140 12152 9168 12180
rect 9324 12152 9352 12192
rect 9481 12189 9493 12192
rect 9527 12189 9539 12223
rect 9481 12183 9539 12189
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9140 12124 9352 12152
rect 9692 12152 9720 12183
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9858 12180 9864 12232
rect 9916 12180 9922 12232
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12222 10839 12223
rect 10870 12222 10876 12232
rect 10827 12194 10876 12222
rect 10827 12189 10839 12194
rect 10781 12183 10839 12189
rect 10870 12180 10876 12194
rect 10928 12180 10934 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11256 12229 11284 12260
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 11624 12220 11652 12260
rect 12713 12233 12771 12239
rect 11701 12223 11759 12229
rect 11701 12220 11713 12223
rect 11624 12192 11713 12220
rect 11701 12189 11713 12192
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 11882 12220 11888 12232
rect 11839 12192 11888 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 10244 12152 10272 12180
rect 9692 12124 10272 12152
rect 10965 12155 11023 12161
rect 10965 12121 10977 12155
rect 11011 12152 11023 12155
rect 11164 12152 11192 12180
rect 11011 12124 11192 12152
rect 11011 12121 11023 12124
rect 10965 12115 11023 12121
rect 11422 12112 11428 12164
rect 11480 12112 11486 12164
rect 12176 12152 12204 12183
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12713 12199 12725 12233
rect 12759 12199 12771 12233
rect 12912 12229 12940 12396
rect 12713 12193 12771 12199
rect 12897 12223 12955 12229
rect 12728 12164 12756 12193
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12345 12155 12403 12161
rect 11541 12124 12296 12152
rect 7006 12084 7012 12096
rect 6840 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9858 12084 9864 12096
rect 9447 12056 9864 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 10413 12087 10471 12093
rect 10413 12053 10425 12087
rect 10459 12084 10471 12087
rect 10502 12084 10508 12096
rect 10459 12056 10508 12084
rect 10459 12053 10471 12056
rect 10413 12047 10471 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 11541 12084 11569 12124
rect 12268 12096 12296 12124
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 12391 12124 12572 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 10928 12056 11569 12084
rect 10928 12044 10934 12056
rect 12250 12044 12256 12096
rect 12308 12044 12314 12096
rect 12434 12044 12440 12096
rect 12492 12093 12498 12096
rect 12492 12047 12501 12093
rect 12544 12084 12572 12124
rect 12710 12112 12716 12164
rect 12768 12112 12774 12164
rect 12802 12084 12808 12096
rect 12544 12056 12808 12084
rect 12492 12044 12498 12047
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 1104 11994 14076 12016
rect 1104 11942 4918 11994
rect 4970 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 5238 11994
rect 5290 11942 10918 11994
rect 10970 11942 10982 11994
rect 11034 11942 11046 11994
rect 11098 11942 11110 11994
rect 11162 11942 11174 11994
rect 11226 11942 11238 11994
rect 11290 11942 14076 11994
rect 1104 11920 14076 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3513 11883 3571 11889
rect 3513 11849 3525 11883
rect 3559 11880 3571 11883
rect 3602 11880 3608 11892
rect 3559 11852 3608 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4522 11840 4528 11892
rect 4580 11840 4586 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7558 11880 7564 11892
rect 7147 11852 7564 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7650 11840 7656 11892
rect 7708 11840 7714 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7760 11852 7849 11880
rect 5810 11812 5816 11824
rect 4632 11784 5816 11812
rect 4632 11756 4660 11784
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3068 11716 3341 11744
rect 3068 11688 3096 11716
rect 3329 11713 3341 11716
rect 3375 11744 3387 11747
rect 4062 11744 4068 11756
rect 3375 11716 4068 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4614 11704 4620 11756
rect 4672 11704 4678 11756
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4890 11744 4896 11756
rect 4755 11716 4896 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 5000 11753 5028 11784
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 7668 11812 7696 11840
rect 7576 11784 7696 11812
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 6362 11744 6368 11756
rect 5215 11716 6368 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7064 11716 7297 11744
rect 7064 11704 7070 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 7576 11753 7604 11784
rect 7760 11753 7788 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 7837 11843 7895 11849
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 7984 11852 9720 11880
rect 7984 11840 7990 11852
rect 9692 11753 9720 11852
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9824 11852 9965 11880
rect 9824 11840 9830 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10229 11883 10287 11889
rect 10100 11852 10180 11880
rect 10100 11840 10106 11852
rect 9858 11772 9864 11824
rect 9916 11772 9922 11824
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 9766 11744 9772 11756
rect 9723 11716 9772 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 3050 11636 3056 11688
rect 3108 11636 3114 11688
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3252 11540 3280 11639
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 3878 11676 3884 11688
rect 3743 11648 3884 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7156 11648 7481 11676
rect 7156 11636 7162 11648
rect 7469 11645 7481 11648
rect 7515 11676 7527 11679
rect 7852 11676 7880 11707
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 9876 11742 9904 11772
rect 10152 11756 10180 11852
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 11514 11880 11520 11892
rect 10275 11852 11520 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11606 11840 11612 11892
rect 11664 11840 11670 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12342 11880 12348 11892
rect 12115 11852 12348 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12434 11840 12440 11892
rect 12492 11840 12498 11892
rect 10042 11742 10048 11756
rect 9876 11714 10048 11742
rect 10042 11704 10048 11714
rect 10100 11704 10106 11756
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10192 11716 10241 11744
rect 10192 11704 10198 11716
rect 10229 11713 10241 11716
rect 10275 11744 10287 11747
rect 10686 11744 10692 11756
rect 10275 11716 10692 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 11624 11744 11652 11840
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11624 11716 11897 11744
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 12452 11753 12480 11840
rect 12428 11747 12486 11753
rect 12428 11713 12440 11747
rect 12474 11713 12486 11747
rect 12428 11707 12486 11713
rect 7515 11648 7880 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 8110 11636 8116 11688
rect 8168 11636 8174 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10410 11676 10416 11688
rect 9999 11648 10416 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 10778 11676 10784 11688
rect 10560 11648 10784 11676
rect 10560 11636 10566 11648
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 11698 11636 11704 11688
rect 11756 11636 11762 11688
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11992 11676 12020 11704
rect 11839 11648 12020 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 7929 11611 7987 11617
rect 7929 11577 7941 11611
rect 7975 11577 7987 11611
rect 8128 11608 8156 11636
rect 10594 11608 10600 11620
rect 8128 11580 10600 11608
rect 7929 11571 7987 11577
rect 4706 11540 4712 11552
rect 3016 11512 4712 11540
rect 3016 11500 3022 11512
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 7944 11540 7972 11571
rect 10594 11568 10600 11580
rect 10652 11568 10658 11620
rect 7432 11512 7972 11540
rect 9769 11543 9827 11549
rect 7432 11500 7438 11512
rect 9769 11509 9781 11543
rect 9815 11540 9827 11543
rect 11330 11540 11336 11552
rect 9815 11512 11336 11540
rect 9815 11509 9827 11512
rect 9769 11503 9827 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 13170 11540 13176 11552
rect 11756 11512 13176 11540
rect 11756 11500 11762 11512
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13538 11500 13544 11552
rect 13596 11500 13602 11552
rect 1104 11450 14076 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 14076 11450
rect 1104 11376 14076 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 2498 11336 2504 11348
rect 1535 11308 2504 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 2498 11296 2504 11308
rect 2556 11336 2562 11348
rect 2556 11308 3648 11336
rect 2556 11296 2562 11308
rect 2866 11160 2872 11212
rect 2924 11160 2930 11212
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3326 11132 3332 11144
rect 3191 11104 3332 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 3620 11141 3648 11308
rect 4246 11296 4252 11348
rect 4304 11296 4310 11348
rect 7374 11296 7380 11348
rect 7432 11296 7438 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11790 11336 11796 11348
rect 11379 11308 11796 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4264 11200 4292 11296
rect 5350 11228 5356 11280
rect 5408 11268 5414 11280
rect 7926 11268 7932 11280
rect 5408 11240 7932 11268
rect 5408 11228 5414 11240
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 10152 11268 10180 11299
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12492 11308 12817 11336
rect 12492 11296 12498 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 12805 11299 12863 11305
rect 13170 11296 13176 11348
rect 13228 11296 13234 11348
rect 10226 11268 10232 11280
rect 9646 11240 10232 11268
rect 3752 11172 4384 11200
rect 3752 11160 3758 11172
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 4246 11132 4252 11144
rect 3651 11104 4252 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4356 11141 4384 11172
rect 4816 11172 6776 11200
rect 4816 11144 4844 11172
rect 6748 11144 6776 11172
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 9646 11200 9674 11240
rect 10226 11228 10232 11240
rect 10284 11268 10290 11280
rect 12342 11268 12348 11280
rect 10284 11240 12348 11268
rect 10284 11228 10290 11240
rect 9456 11172 9674 11200
rect 9456 11160 9462 11172
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10873 11203 10931 11209
rect 10008 11172 10088 11200
rect 10008 11160 10014 11172
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 4890 11092 4896 11144
rect 4948 11132 4954 11144
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4948 11104 4997 11132
rect 4948 11092 4954 11104
rect 4985 11101 4997 11104
rect 5031 11132 5043 11135
rect 5810 11132 5816 11144
rect 5031 11104 5816 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 2624 11067 2682 11073
rect 2624 11033 2636 11067
rect 2670 11064 2682 11067
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2670 11036 2973 11064
rect 2670 11033 2682 11036
rect 2624 11027 2682 11033
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 4764 11036 5948 11064
rect 4764 11024 4770 11036
rect 5920 11008 5948 11036
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 6472 11064 6500 11095
rect 6420 11036 6500 11064
rect 6656 11064 6684 11095
rect 6730 11092 6736 11144
rect 6788 11092 6794 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 10060 11141 10088 11172
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 10919 11172 11437 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7340 11104 7389 11132
rect 7340 11092 7346 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 10045 11135 10103 11141
rect 7377 11095 7435 11101
rect 8496 11104 9996 11132
rect 7300 11064 7328 11092
rect 8496 11076 8524 11104
rect 8294 11064 8300 11076
rect 6656 11036 7328 11064
rect 7383 11036 8300 11064
rect 6420 11024 6426 11036
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4893 10999 4951 11005
rect 4893 10996 4905 10999
rect 4580 10968 4905 10996
rect 4580 10956 4586 10968
rect 4893 10965 4905 10968
rect 4939 10965 4951 10999
rect 4893 10959 4951 10965
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6549 10999 6607 11005
rect 6549 10996 6561 10999
rect 6052 10968 6561 10996
rect 6052 10956 6058 10968
rect 6549 10965 6561 10968
rect 6595 10996 6607 10999
rect 7383 10996 7411 11036
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 8478 11024 8484 11076
rect 8536 11024 8542 11076
rect 9968 11064 9996 11104
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 10778 11132 10784 11144
rect 10459 11104 10784 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11330 11132 11336 11144
rect 11195 11104 11336 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11716 11141 11744 11240
rect 12342 11228 12348 11240
rect 12400 11268 12406 11280
rect 13538 11268 13544 11280
rect 12400 11240 13544 11268
rect 12400 11228 12406 11240
rect 11808 11172 12848 11200
rect 11808 11141 11836 11172
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11422 11064 11428 11076
rect 9692 11036 9904 11064
rect 9968 11036 11428 11064
rect 6595 10968 7411 10996
rect 6595 10965 6607 10968
rect 6549 10959 6607 10965
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9692 10996 9720 11036
rect 9876 11008 9904 11036
rect 11422 11024 11428 11036
rect 11480 11064 11486 11076
rect 11808 11064 11836 11095
rect 11480 11036 11836 11064
rect 11900 11064 11928 11095
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12360 11141 12388 11172
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12176 11064 12204 11095
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12820 11141 12848 11172
rect 12912 11144 12940 11240
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12894 11092 12900 11144
rect 12952 11092 12958 11144
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 11900 11036 12204 11064
rect 12360 11036 12449 11064
rect 11480 11024 11486 11036
rect 11900 11008 11928 11036
rect 12360 11008 12388 11036
rect 12437 11033 12449 11036
rect 12483 11033 12495 11067
rect 12437 11027 12495 11033
rect 9364 10968 9720 10996
rect 9364 10956 9370 10968
rect 9766 10956 9772 11008
rect 9824 10956 9830 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 9916 10968 10333 10996
rect 9916 10956 9922 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 11054 10996 11060 11008
rect 10744 10968 11060 10996
rect 10744 10956 10750 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 11882 10956 11888 11008
rect 11940 10956 11946 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12584 10968 12725 10996
rect 12584 10956 12590 10968
rect 12713 10965 12725 10968
rect 12759 10965 12771 10999
rect 12713 10959 12771 10965
rect 1104 10906 14076 10928
rect 1104 10854 4918 10906
rect 4970 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 5238 10906
rect 5290 10854 10918 10906
rect 10970 10854 10982 10906
rect 11034 10854 11046 10906
rect 11098 10854 11110 10906
rect 11162 10854 11174 10906
rect 11226 10854 11238 10906
rect 11290 10854 14076 10906
rect 1104 10832 14076 10854
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3476 10764 3525 10792
rect 3476 10752 3482 10764
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 3936 10764 4721 10792
rect 3936 10752 3942 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 5994 10792 6000 10804
rect 4709 10755 4767 10761
rect 4908 10764 6000 10792
rect 3068 10696 3740 10724
rect 3068 10600 3096 10696
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3712 10665 3740 10696
rect 4522 10684 4528 10736
rect 4580 10684 4586 10736
rect 3697 10659 3755 10665
rect 3384 10628 3464 10656
rect 3384 10616 3390 10628
rect 2958 10548 2964 10600
rect 3016 10548 3022 10600
rect 3050 10548 3056 10600
rect 3108 10548 3114 10600
rect 3436 10597 3464 10628
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3697 10619 3755 10625
rect 3804 10628 3985 10656
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3602 10588 3608 10600
rect 3421 10551 3479 10557
rect 3528 10560 3608 10588
rect 3251 10520 3279 10551
rect 3528 10520 3556 10560
rect 3602 10548 3608 10560
rect 3660 10588 3666 10600
rect 3804 10588 3832 10628
rect 3973 10625 3985 10628
rect 4019 10656 4031 10659
rect 4062 10656 4068 10668
rect 4019 10628 4068 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4540 10656 4568 10684
rect 4908 10665 4936 10764
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7432 10764 7573 10792
rect 7432 10752 7438 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 8386 10792 8392 10804
rect 7699 10764 8392 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9180 10764 9628 10792
rect 9180 10752 9186 10764
rect 5184 10696 5488 10724
rect 5184 10665 5212 10696
rect 4212 10628 4568 10656
rect 4893 10659 4951 10665
rect 4212 10616 4218 10628
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5316 10628 5365 10656
rect 5316 10616 5322 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5460 10656 5488 10696
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 6788 10696 7420 10724
rect 6788 10684 6794 10696
rect 5534 10656 5540 10668
rect 5460 10628 5540 10656
rect 5353 10619 5411 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 3660 10560 3832 10588
rect 3881 10591 3939 10597
rect 3660 10548 3666 10560
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 5626 10588 5632 10600
rect 3927 10560 5632 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 3251 10492 3556 10520
rect 3786 10480 3792 10532
rect 3844 10480 3850 10532
rect 4798 10480 4804 10532
rect 4856 10520 4862 10532
rect 4985 10523 5043 10529
rect 4985 10520 4997 10523
rect 4856 10492 4997 10520
rect 4856 10480 4862 10492
rect 4985 10489 4997 10492
rect 5031 10489 5043 10523
rect 4985 10483 5043 10489
rect 5077 10523 5135 10529
rect 5077 10489 5089 10523
rect 5123 10489 5135 10523
rect 5828 10520 5856 10619
rect 6362 10616 6368 10668
rect 6420 10654 6426 10668
rect 6457 10659 6515 10665
rect 6457 10654 6469 10659
rect 6420 10626 6469 10654
rect 6420 10616 6426 10626
rect 6457 10625 6469 10626
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6696 10628 6929 10656
rect 6696 10616 6702 10628
rect 6917 10625 6929 10628
rect 6963 10656 6975 10659
rect 7282 10656 7288 10668
rect 6963 10628 7288 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7392 10665 7420 10696
rect 8036 10696 8524 10724
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7616 10628 7757 10656
rect 7616 10616 7622 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8036 10665 8064 10696
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7892 10628 7941 10656
rect 7892 10616 7898 10628
rect 7929 10625 7941 10628
rect 7975 10656 7987 10659
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7975 10628 8033 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 5951 10560 6561 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6549 10557 6561 10560
rect 6595 10588 6607 10591
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6595 10560 6745 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 6733 10557 6745 10560
rect 6779 10588 6791 10591
rect 7190 10588 7196 10600
rect 6779 10560 7196 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 7190 10548 7196 10560
rect 7248 10588 7254 10600
rect 7650 10588 7656 10600
rect 7248 10560 7656 10588
rect 7248 10548 7254 10560
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8110 10548 8116 10600
rect 8168 10548 8174 10600
rect 8220 10588 8248 10619
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8496 10665 8524 10696
rect 9600 10668 9628 10764
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9732 10764 9781 10792
rect 9732 10752 9738 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 9858 10752 9864 10804
rect 9916 10752 9922 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10134 10792 10140 10804
rect 10008 10764 10140 10792
rect 10008 10752 10014 10764
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10376 10764 10517 10792
rect 10376 10752 10382 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 10686 10752 10692 10804
rect 10744 10752 10750 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11330 10792 11336 10804
rect 11103 10764 11336 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11514 10752 11520 10804
rect 11572 10752 11578 10804
rect 11606 10752 11612 10804
rect 11664 10752 11670 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12253 10795 12311 10801
rect 12253 10792 12265 10795
rect 12032 10764 12265 10792
rect 12032 10752 12038 10764
rect 12253 10761 12265 10764
rect 12299 10761 12311 10795
rect 12253 10755 12311 10761
rect 12618 10752 12624 10804
rect 12676 10752 12682 10804
rect 10410 10724 10416 10736
rect 9692 10696 10416 10724
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8527 10628 9137 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 8570 10588 8576 10600
rect 8220 10560 8576 10588
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 9232 10588 9260 10619
rect 9582 10616 9588 10668
rect 9640 10616 9646 10668
rect 9692 10665 9720 10696
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 10704 10724 10732 10752
rect 11238 10724 11244 10736
rect 10704 10696 11244 10724
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9950 10656 9956 10668
rect 9677 10619 9735 10625
rect 9876 10628 9956 10656
rect 9876 10588 9904 10628
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 10100 10628 10149 10656
rect 10100 10616 10106 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10836 10628 10885 10656
rect 10836 10616 10842 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 11532 10656 11560 10752
rect 11624 10724 11652 10752
rect 12805 10727 12863 10733
rect 12805 10724 12817 10727
rect 11624 10696 12817 10724
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11532 10628 11713 10656
rect 10873 10619 10931 10625
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 12066 10656 12072 10668
rect 11701 10619 11759 10625
rect 11808 10628 12072 10656
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9232 10560 9904 10588
rect 9968 10560 10241 10588
rect 6086 10520 6092 10532
rect 5828 10492 6092 10520
rect 5077 10483 5135 10489
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5092 10452 5120 10483
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 6178 10480 6184 10532
rect 6236 10480 6242 10532
rect 6362 10480 6368 10532
rect 6420 10520 6426 10532
rect 6420 10492 7604 10520
rect 6420 10480 6426 10492
rect 7208 10464 7236 10492
rect 4580 10424 5120 10452
rect 4580 10412 4586 10424
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5813 10455 5871 10461
rect 5813 10452 5825 10455
rect 5500 10424 5825 10452
rect 5500 10412 5506 10424
rect 5813 10421 5825 10424
rect 5859 10452 5871 10455
rect 6454 10452 6460 10464
rect 5859 10424 6460 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 7098 10452 7104 10464
rect 6604 10424 7104 10452
rect 6604 10412 6610 10424
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7190 10412 7196 10464
rect 7248 10412 7254 10464
rect 7576 10452 7604 10492
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 7800 10492 9505 10520
rect 7800 10480 7806 10492
rect 9493 10489 9505 10492
rect 9539 10489 9551 10523
rect 9968 10520 9996 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 10502 10588 10508 10600
rect 10275 10560 10508 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10888 10588 10916 10619
rect 11808 10588 11836 10628
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12360 10665 12388 10696
rect 12805 10693 12817 10696
rect 12851 10693 12863 10727
rect 12805 10687 12863 10693
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 10888 10560 11836 10588
rect 11974 10548 11980 10600
rect 12032 10548 12038 10600
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 12526 10588 12532 10600
rect 12483 10560 12532 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 12894 10588 12900 10600
rect 12667 10560 12900 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 9493 10483 9551 10489
rect 9692 10492 9996 10520
rect 9692 10464 9720 10492
rect 10042 10480 10048 10532
rect 10100 10480 10106 10532
rect 12636 10520 12664 10551
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 12452 10492 12664 10520
rect 12452 10464 12480 10492
rect 9214 10452 9220 10464
rect 7576 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9674 10412 9680 10464
rect 9732 10412 9738 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 9916 10424 10149 10452
rect 9916 10412 9922 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 11790 10412 11796 10464
rect 11848 10412 11854 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 1104 10362 14076 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 14076 10362
rect 1104 10288 14076 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 4801 10251 4859 10257
rect 4801 10248 4813 10251
rect 2924 10220 4813 10248
rect 2924 10208 2930 10220
rect 4801 10217 4813 10220
rect 4847 10217 4859 10251
rect 4801 10211 4859 10217
rect 6178 10208 6184 10260
rect 6236 10208 6242 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7340 10220 8984 10248
rect 7340 10208 7346 10220
rect 3418 10072 3424 10124
rect 3476 10072 3482 10124
rect 6196 10112 6224 10208
rect 8386 10180 8392 10192
rect 7944 10152 8392 10180
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6196 10084 6929 10112
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 7944 10121 7972 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7432 10084 7573 10112
rect 7432 10072 7438 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8110 10072 8116 10124
rect 8168 10072 8174 10124
rect 8404 10112 8432 10140
rect 8570 10112 8576 10124
rect 8404 10084 8576 10112
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3252 9976 3280 10007
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10044 4307 10047
rect 6546 10044 6552 10056
rect 4295 10016 6552 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10013 7067 10047
rect 7009 10007 7067 10013
rect 3252 9948 3372 9976
rect 3344 9920 3372 9948
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 4338 9976 4344 9988
rect 3936 9948 4344 9976
rect 3936 9936 3942 9948
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4614 9976 4620 9988
rect 4479 9948 4620 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 6822 9976 6828 9988
rect 6319 9948 6828 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 7024 9920 7052 10007
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7484 9976 7512 10007
rect 7650 10004 7656 10056
rect 7708 10053 7714 10056
rect 7708 10047 7757 10053
rect 7708 10013 7711 10047
rect 7745 10013 7757 10047
rect 7708 10007 7757 10013
rect 7708 10004 7714 10007
rect 7834 10004 7840 10056
rect 7892 10044 7898 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7892 10016 8033 10044
rect 7892 10004 7898 10016
rect 8021 10013 8033 10016
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8956 10053 8984 10220
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 12158 10208 12164 10260
rect 12216 10208 12222 10260
rect 9950 10180 9956 10192
rect 9784 10152 9956 10180
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8352 10016 8401 10044
rect 8352 10004 8358 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 8389 10007 8447 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9030 10004 9036 10056
rect 9088 10004 9094 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9214 10044 9220 10056
rect 9171 10016 9220 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9784 10053 9812 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 12802 10180 12808 10192
rect 11480 10152 12808 10180
rect 11480 10140 11486 10152
rect 12802 10140 12808 10152
rect 12860 10140 12866 10192
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9968 10084 10333 10112
rect 9968 10056 9996 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 9048 9976 9076 10004
rect 7484 9948 9076 9976
rect 9508 9976 9536 10007
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 9950 10004 9956 10056
rect 10008 10004 10014 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10134 10044 10140 10056
rect 10091 10016 10140 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10336 10016 10824 10044
rect 10336 9976 10364 10016
rect 10796 9988 10824 10016
rect 9508 9948 10364 9976
rect 10413 9979 10471 9985
rect 10413 9945 10425 9979
rect 10459 9945 10471 9979
rect 10413 9939 10471 9945
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2924 9880 2973 9908
rect 2924 9868 2930 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 3326 9868 3332 9920
rect 3384 9868 3390 9920
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3660 9880 4077 9908
rect 3660 9868 3666 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 4212 9880 6469 9908
rect 4212 9868 4218 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 7006 9868 7012 9920
rect 7064 9868 7070 9920
rect 7282 9868 7288 9920
rect 7340 9868 7346 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7616 9880 7849 9908
rect 7616 9868 7622 9880
rect 7837 9877 7849 9880
rect 7883 9908 7895 9911
rect 8386 9908 8392 9920
rect 7883 9880 8392 9908
rect 7883 9877 7895 9880
rect 7837 9871 7895 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8536 9880 9045 9908
rect 8536 9868 8542 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 9214 9868 9220 9920
rect 9272 9868 9278 9920
rect 10428 9908 10456 9939
rect 10502 9936 10508 9988
rect 10560 9976 10566 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10560 9948 10701 9976
rect 10560 9936 10566 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 10778 9936 10784 9988
rect 10836 9936 10842 9988
rect 10594 9908 10600 9920
rect 10428 9880 10600 9908
rect 10594 9868 10600 9880
rect 10652 9908 10658 9920
rect 11790 9908 11796 9920
rect 10652 9880 11796 9908
rect 10652 9868 10658 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 1104 9818 14076 9840
rect 1104 9766 4918 9818
rect 4970 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 5238 9818
rect 5290 9766 10918 9818
rect 10970 9766 10982 9818
rect 11034 9766 11046 9818
rect 11098 9766 11110 9818
rect 11162 9766 11174 9818
rect 11226 9766 11238 9818
rect 11290 9766 14076 9818
rect 1104 9744 14076 9766
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3970 9704 3976 9716
rect 3292 9676 3976 9704
rect 3292 9664 3298 9676
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 4157 9707 4215 9713
rect 4157 9674 4169 9707
rect 4080 9673 4169 9674
rect 4203 9673 4215 9707
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4080 9667 4215 9673
rect 4264 9676 4629 9704
rect 4080 9646 4200 9667
rect 4080 9636 4108 9646
rect 4007 9608 4108 9636
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2087 9540 2176 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2148 9509 2176 9540
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3292 9540 3433 9568
rect 3292 9528 3298 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 4007 9568 4035 9608
rect 4264 9568 4292 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 5810 9704 5816 9716
rect 4617 9667 4675 9673
rect 5000 9676 5816 9704
rect 4890 9596 4896 9648
rect 4948 9596 4954 9648
rect 3421 9531 3479 9537
rect 3528 9540 4035 9568
rect 4080 9540 4292 9568
rect 4341 9574 4399 9577
rect 4522 9574 4528 9580
rect 4341 9571 4528 9574
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 2639 9472 2789 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2958 9460 2964 9512
rect 3016 9460 3022 9512
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 2317 9435 2375 9441
rect 2317 9401 2329 9435
rect 2363 9432 2375 9435
rect 2866 9432 2872 9444
rect 2363 9404 2872 9432
rect 2363 9401 2375 9404
rect 2317 9395 2375 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1820 9336 1869 9364
rect 1820 9324 1826 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 3252 9364 3280 9528
rect 3528 9512 3556 9540
rect 3326 9460 3332 9512
rect 3384 9460 3390 9512
rect 3510 9460 3516 9512
rect 3568 9460 3574 9512
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4080 9509 4108 9540
rect 4341 9537 4353 9571
rect 4387 9546 4528 9571
rect 4387 9537 4399 9546
rect 4341 9531 4399 9537
rect 4522 9528 4528 9546
rect 4580 9528 4586 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4706 9568 4712 9580
rect 4663 9540 4712 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4908 9568 4936 9596
rect 5000 9577 5028 9676
rect 5810 9664 5816 9676
rect 5868 9704 5874 9716
rect 7282 9704 7288 9716
rect 5868 9676 7288 9704
rect 5868 9664 5874 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 8386 9704 8392 9716
rect 8220 9676 8392 9704
rect 6086 9636 6092 9648
rect 5920 9608 6092 9636
rect 4816 9540 4936 9568
rect 4985 9571 5043 9577
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4246 9500 4252 9512
rect 4111 9472 4252 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4816 9500 4844 9540
rect 4985 9537 4997 9571
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5626 9568 5632 9580
rect 5399 9540 5632 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 5920 9577 5948 9608
rect 6086 9596 6092 9608
rect 6144 9636 6150 9648
rect 7006 9636 7012 9648
rect 6144 9608 7012 9636
rect 6144 9596 6150 9608
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 8220 9636 8248 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8481 9707 8539 9713
rect 8481 9673 8493 9707
rect 8527 9673 8539 9707
rect 8481 9667 8539 9673
rect 8496 9636 8524 9667
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 9033 9707 9091 9713
rect 9033 9704 9045 9707
rect 8628 9676 9045 9704
rect 8628 9664 8634 9676
rect 9033 9673 9045 9676
rect 9079 9673 9091 9707
rect 9033 9667 9091 9673
rect 10318 9664 10324 9716
rect 10376 9664 10382 9716
rect 10870 9704 10876 9716
rect 10796 9676 10876 9704
rect 8662 9636 8668 9648
rect 8220 9608 8285 9636
rect 8496 9608 8668 9636
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6730 9568 6736 9580
rect 6227 9540 6736 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 4479 9472 4844 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 6012 9500 6040 9531
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7024 9540 7205 9568
rect 6638 9500 6644 9512
rect 4948 9472 6644 9500
rect 4948 9460 4954 9472
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 3344 9432 3372 9460
rect 5537 9435 5595 9441
rect 5537 9432 5549 9435
rect 3344 9404 5549 9432
rect 5537 9401 5549 9404
rect 5583 9401 5595 9435
rect 5537 9395 5595 9401
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 6748 9432 6776 9528
rect 7024 9512 7052 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 5684 9404 6776 9432
rect 5684 9392 5690 9404
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 7300 9432 7328 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 8257 9577 8285 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 9214 9636 9220 9648
rect 8864 9608 9220 9636
rect 8864 9580 8892 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 10336 9636 10364 9664
rect 10796 9636 10824 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 12066 9704 12072 9716
rect 11716 9676 12072 9704
rect 10336 9608 10824 9636
rect 8242 9571 8300 9577
rect 8242 9537 8254 9571
rect 8288 9537 8300 9571
rect 8242 9531 8300 9537
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9568 8447 9571
rect 8478 9568 8484 9580
rect 8435 9540 8484 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9582 9568 9588 9580
rect 9171 9540 9588 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8110 9500 8116 9512
rect 8067 9472 8116 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 9140 9500 9168 9531
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10100 9540 10149 9568
rect 10100 9528 10106 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 10796 9577 10824 9608
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 11716 9645 11744 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 11388 9608 11529 9636
rect 11388 9596 11394 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 11517 9599 11575 9605
rect 11701 9639 11759 9645
rect 11701 9605 11713 9639
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 11885 9639 11943 9645
rect 11885 9605 11897 9639
rect 11931 9636 11943 9639
rect 12434 9636 12440 9648
rect 11931 9608 12440 9636
rect 11931 9605 11943 9608
rect 11885 9599 11943 9605
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10468 9540 10517 9568
rect 10468 9528 10474 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9537 10655 9571
rect 10597 9531 10655 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 8812 9472 9168 9500
rect 10244 9500 10272 9528
rect 10612 9500 10640 9531
rect 10244 9472 10640 9500
rect 8812 9460 8818 9472
rect 6880 9404 7328 9432
rect 6880 9392 6886 9404
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 8628 9404 9873 9432
rect 8628 9392 8634 9404
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 9861 9395 9919 9401
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 3252 9336 6929 9364
rect 1857 9327 1915 9333
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7745 9367 7803 9373
rect 7745 9364 7757 9367
rect 7156 9336 7757 9364
rect 7156 9324 7162 9336
rect 7745 9333 7757 9336
rect 7791 9333 7803 9367
rect 7745 9327 7803 9333
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 8168 9336 8677 9364
rect 8168 9324 8174 9336
rect 8665 9333 8677 9336
rect 8711 9364 8723 9367
rect 8938 9364 8944 9376
rect 8711 9336 8944 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 8938 9324 8944 9336
rect 8996 9364 9002 9376
rect 9674 9364 9680 9376
rect 8996 9336 9680 9364
rect 8996 9324 9002 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10888 9364 10916 9531
rect 10962 9528 10968 9580
rect 11020 9558 11026 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11020 9530 11055 9558
rect 11164 9540 11989 9568
rect 11020 9528 11026 9530
rect 10966 9527 10978 9528
rect 11012 9527 11024 9528
rect 10966 9521 11024 9527
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 11164 9432 11192 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 12176 9500 12204 9531
rect 11572 9472 12204 9500
rect 11572 9460 11578 9472
rect 11020 9404 11192 9432
rect 11241 9435 11299 9441
rect 11020 9392 11026 9404
rect 11241 9401 11253 9435
rect 11287 9432 11299 9435
rect 12710 9432 12716 9444
rect 11287 9404 12716 9432
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 10744 9336 10916 9364
rect 10744 9324 10750 9336
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11756 9336 11989 9364
rect 11756 9324 11762 9336
rect 11977 9333 11989 9336
rect 12023 9364 12035 9367
rect 12342 9364 12348 9376
rect 12023 9336 12348 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 1104 9274 14076 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 14076 9274
rect 1104 9200 14076 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3418 9160 3424 9172
rect 2915 9132 3424 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3418 9120 3424 9132
rect 3476 9160 3482 9172
rect 4062 9160 4068 9172
rect 3476 9132 4068 9160
rect 3476 9120 3482 9132
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4396 9132 4568 9160
rect 4396 9120 4402 9132
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3436 9064 3893 9092
rect 3436 9036 3464 9064
rect 3881 9061 3893 9064
rect 3927 9061 3939 9095
rect 4430 9092 4436 9104
rect 3881 9055 3939 9061
rect 4080 9064 4436 9092
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3016 8996 3157 9024
rect 3016 8984 3022 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 3418 8984 3424 9036
rect 3476 8984 3482 9036
rect 3602 8984 3608 9036
rect 3660 8984 3666 9036
rect 4080 9033 4108 9064
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 4540 9092 4568 9132
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 4856 9132 5365 9160
rect 4856 9120 4862 9132
rect 4890 9092 4896 9104
rect 4540 9064 4896 9092
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4246 9024 4252 9036
rect 4065 8987 4123 8993
rect 4172 8996 4252 9024
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8956 1547 8959
rect 2774 8956 2780 8968
rect 1535 8928 2780 8956
rect 1535 8925 1547 8928
rect 1489 8919 1547 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3108 8928 3249 8956
rect 3108 8916 3114 8928
rect 3237 8925 3249 8928
rect 3283 8956 3295 8959
rect 3970 8956 3976 8968
rect 3283 8928 3976 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4172 8965 4200 8996
rect 4246 8984 4252 8996
rect 4304 9024 4310 9036
rect 4304 8996 4660 9024
rect 4304 8984 4310 8996
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 1762 8897 1768 8900
rect 1756 8888 1768 8897
rect 1723 8860 1768 8888
rect 1756 8851 1768 8860
rect 1762 8848 1768 8851
rect 1820 8848 1826 8900
rect 4172 8888 4200 8919
rect 4338 8916 4344 8968
rect 4396 8916 4402 8968
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 4632 8965 4660 8996
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 4764 8996 4844 9024
rect 4764 8984 4770 8996
rect 4816 8965 4844 8996
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 3436 8860 4200 8888
rect 2958 8780 2964 8832
rect 3016 8780 3022 8832
rect 3436 8829 3464 8860
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 4356 8829 4384 8916
rect 4632 8888 4660 8919
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 5005 8959 5063 8965
rect 5005 8958 5017 8959
rect 5000 8928 5017 8958
rect 5005 8925 5017 8928
rect 5051 8958 5063 8959
rect 5184 8958 5212 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 5592 9132 6377 9160
rect 5592 9120 5598 9132
rect 6365 9129 6377 9132
rect 6411 9129 6423 9163
rect 6365 9123 6423 9129
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 7098 9160 7104 9172
rect 6696 9132 7104 9160
rect 6696 9120 6702 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 7432 9132 7573 9160
rect 7432 9120 7438 9132
rect 7561 9129 7573 9132
rect 7607 9129 7619 9163
rect 7561 9123 7619 9129
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8938 9160 8944 9172
rect 7975 9132 8944 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5626 9092 5632 9104
rect 5307 9064 5632 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 7650 9092 7656 9104
rect 6564 9064 7656 9092
rect 5810 9024 5816 9036
rect 5736 8996 5816 9024
rect 5051 8930 5212 8958
rect 5051 8925 5063 8930
rect 5005 8919 5063 8925
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5736 8965 5764 8996
rect 5810 8984 5816 8996
rect 5868 9024 5874 9036
rect 6362 9024 6368 9036
rect 5868 8996 6368 9024
rect 5868 8984 5874 8996
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5500 8928 5549 8956
rect 5500 8916 5506 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6564 8965 6592 9064
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 7006 9024 7012 9036
rect 6932 8996 7012 9024
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 6932 8965 6960 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7944 9024 7972 9123
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9030 9120 9036 9172
rect 9088 9120 9094 9172
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 10410 9120 10416 9172
rect 10468 9120 10474 9172
rect 10962 9120 10968 9172
rect 11020 9120 11026 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11514 9160 11520 9172
rect 11112 9132 11520 9160
rect 11112 9120 11118 9132
rect 11514 9120 11520 9132
rect 11572 9160 11578 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11572 9132 11897 9160
rect 11572 9120 11578 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 8846 9052 8852 9104
rect 8904 9052 8910 9104
rect 9309 9095 9367 9101
rect 9309 9061 9321 9095
rect 9355 9092 9367 9095
rect 9674 9092 9680 9104
rect 9355 9064 9680 9092
rect 9355 9061 9367 9064
rect 9309 9055 9367 9061
rect 9674 9052 9680 9064
rect 9732 9092 9738 9104
rect 10134 9092 10140 9104
rect 9732 9064 10140 9092
rect 9732 9052 9738 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10336 9092 10364 9120
rect 11241 9095 11299 9101
rect 11241 9092 11253 9095
rect 10336 9064 11253 9092
rect 11241 9061 11253 9064
rect 11287 9061 11299 9095
rect 11241 9055 11299 9061
rect 7300 8996 7972 9024
rect 7300 8968 7328 8996
rect 6926 8959 6984 8965
rect 6926 8925 6938 8959
rect 6972 8925 6984 8959
rect 6926 8919 6984 8925
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 7558 8956 7564 8968
rect 7392 8928 7564 8956
rect 4706 8888 4712 8900
rect 4632 8860 4712 8888
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 6840 8888 6868 8916
rect 6227 8860 6868 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7392 8888 7420 8928
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7708 8928 7757 8956
rect 7708 8916 7714 8928
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7892 8928 7941 8956
rect 7892 8916 7898 8928
rect 7929 8925 7941 8928
rect 7975 8956 7987 8959
rect 8864 8956 8892 9052
rect 10318 9024 10324 9036
rect 8956 8996 10324 9024
rect 8956 8965 8984 8996
rect 10318 8984 10324 8996
rect 10376 9024 10382 9036
rect 10686 9024 10692 9036
rect 10376 8996 10692 9024
rect 10376 8984 10382 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10888 8996 11560 9024
rect 10888 8968 10916 8996
rect 7975 8928 8892 8956
rect 8941 8959 8999 8965
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9306 8956 9312 8968
rect 9263 8928 9312 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 9582 8956 9588 8968
rect 9539 8928 9588 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 9582 8916 9588 8928
rect 9640 8956 9646 8968
rect 10538 8959 10596 8965
rect 10538 8956 10550 8959
rect 9640 8928 10550 8956
rect 9640 8916 9646 8928
rect 10538 8925 10550 8928
rect 10584 8925 10596 8959
rect 10538 8919 10596 8925
rect 10870 8916 10876 8968
rect 10928 8916 10934 8968
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 7156 8860 7420 8888
rect 7469 8891 7527 8897
rect 7156 8848 7162 8860
rect 7469 8857 7481 8891
rect 7515 8888 7527 8891
rect 8386 8888 8392 8900
rect 7515 8860 8392 8888
rect 7515 8857 7527 8860
rect 7469 8851 7527 8857
rect 8386 8848 8392 8860
rect 8444 8888 8450 8900
rect 9858 8888 9864 8900
rect 8444 8860 9864 8888
rect 8444 8848 8450 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 11164 8888 11192 8919
rect 11330 8916 11336 8968
rect 11388 8916 11394 8968
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11532 8965 11560 8996
rect 11624 8996 12020 9024
rect 11624 8965 11652 8996
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11992 8956 12020 8996
rect 12158 8984 12164 9036
rect 12216 8984 12222 9036
rect 12417 8959 12475 8965
rect 12417 8956 12429 8959
rect 11992 8928 12429 8956
rect 11701 8919 11759 8925
rect 12417 8925 12429 8928
rect 12463 8925 12475 8959
rect 12417 8919 12475 8925
rect 10100 8860 11192 8888
rect 11440 8888 11468 8916
rect 11716 8888 11744 8919
rect 11440 8860 11744 8888
rect 10100 8848 10106 8860
rect 11974 8848 11980 8900
rect 12032 8848 12038 8900
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 3568 8792 4353 8820
rect 3568 8780 3574 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4614 8820 4620 8832
rect 4479 8792 4620 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4614 8780 4620 8792
rect 4672 8820 4678 8832
rect 4982 8820 4988 8832
rect 4672 8792 4988 8820
rect 4672 8780 4678 8792
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5500 8792 5825 8820
rect 5500 8780 5506 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 8478 8820 8484 8832
rect 7064 8792 8484 8820
rect 7064 8780 7070 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 10410 8820 10416 8832
rect 10192 8792 10416 8820
rect 10192 8780 10198 8792
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10594 8780 10600 8832
rect 10652 8780 10658 8832
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 1104 8730 14076 8752
rect 1104 8678 4918 8730
rect 4970 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 5238 8730
rect 5290 8678 10918 8730
rect 10970 8678 10982 8730
rect 11034 8678 11046 8730
rect 11098 8678 11110 8730
rect 11162 8678 11174 8730
rect 11226 8678 11238 8730
rect 11290 8678 14076 8730
rect 1104 8656 14076 8678
rect 2958 8576 2964 8628
rect 3016 8576 3022 8628
rect 3786 8576 3792 8628
rect 3844 8576 3850 8628
rect 4246 8576 4252 8628
rect 4304 8576 4310 8628
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4396 8588 4445 8616
rect 4396 8576 4402 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 5442 8616 5448 8628
rect 4580 8588 5448 8616
rect 4580 8576 4586 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 6972 8588 8033 8616
rect 6972 8576 6978 8588
rect 8021 8585 8033 8588
rect 8067 8616 8079 8619
rect 10502 8616 10508 8628
rect 8067 8588 10508 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 2976 8548 3004 8576
rect 3237 8551 3295 8557
rect 3237 8548 3249 8551
rect 2976 8520 3249 8548
rect 3237 8517 3249 8520
rect 3283 8517 3295 8551
rect 3237 8511 3295 8517
rect 3804 8480 3832 8576
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 5828 8548 5856 8576
rect 7282 8548 7288 8560
rect 4120 8520 5856 8548
rect 7208 8520 7288 8548
rect 4120 8508 4126 8520
rect 3252 8452 3832 8480
rect 2961 8347 3019 8353
rect 2961 8313 2973 8347
rect 3007 8344 3019 8347
rect 3252 8344 3280 8452
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 4028 8452 4200 8480
rect 4028 8440 4034 8452
rect 4172 8421 4200 8452
rect 4522 8440 4528 8492
rect 4580 8440 4586 8492
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 7208 8489 7236 8520
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 14182 8548 14188 8560
rect 9355 8520 14188 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10778 8480 10784 8492
rect 10459 8452 10784 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12492 8452 12817 8480
rect 12492 8440 12498 8452
rect 12805 8449 12817 8452
rect 12851 8480 12863 8483
rect 13538 8480 13544 8492
rect 12851 8452 13544 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3881 8415 3939 8421
rect 3881 8412 3893 8415
rect 3375 8384 3893 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3881 8381 3893 8384
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8381 4123 8415
rect 4065 8375 4123 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4203 8384 4752 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 3007 8316 3280 8344
rect 3007 8313 3019 8316
rect 2961 8307 3019 8313
rect 3418 8304 3424 8356
rect 3476 8344 3482 8356
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 3476 8316 3617 8344
rect 3476 8304 3482 8316
rect 3605 8313 3617 8316
rect 3651 8313 3663 8347
rect 3605 8307 3663 8313
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4080 8344 4108 8375
rect 3752 8316 4108 8344
rect 3752 8304 3758 8316
rect 4724 8288 4752 8384
rect 4890 8372 4896 8424
rect 4948 8372 4954 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5902 8412 5908 8424
rect 5123 8384 5908 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5000 8344 5028 8375
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 7650 8412 7656 8424
rect 6420 8384 7656 8412
rect 6420 8372 6426 8384
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 5000 8316 7052 8344
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 3786 8236 3792 8288
rect 3844 8236 3850 8288
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 4706 8236 4712 8288
rect 4764 8236 4770 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5000 8276 5028 8316
rect 7024 8288 7052 8316
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 9122 8344 9128 8356
rect 8444 8316 9128 8344
rect 8444 8304 8450 8316
rect 9122 8304 9128 8316
rect 9180 8344 9186 8356
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 9180 8316 10517 8344
rect 9180 8304 9186 8316
rect 9508 8288 9536 8316
rect 10505 8313 10517 8316
rect 10551 8313 10563 8347
rect 10505 8307 10563 8313
rect 4948 8248 5028 8276
rect 4948 8236 4954 8248
rect 7006 8236 7012 8288
rect 7064 8236 7070 8288
rect 9490 8236 9496 8288
rect 9548 8236 9554 8288
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12621 8279 12679 8285
rect 12621 8276 12633 8279
rect 12216 8248 12633 8276
rect 12216 8236 12222 8248
rect 12621 8245 12633 8248
rect 12667 8245 12679 8279
rect 12621 8239 12679 8245
rect 1104 8186 14076 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 14076 8186
rect 1104 8112 14076 8134
rect 5626 8032 5632 8084
rect 5684 8032 5690 8084
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 6880 8044 7757 8072
rect 6880 8032 6886 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7892 8044 8125 8072
rect 7892 8032 7898 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 10100 8044 10517 8072
rect 10100 8032 10106 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 10652 8044 11529 8072
rect 10652 8032 10658 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 11517 8035 11575 8041
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12032 8044 12265 8072
rect 12032 8032 12038 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8041 12495 8075
rect 12437 8035 12495 8041
rect 5644 7936 5672 8032
rect 11241 8007 11299 8013
rect 11241 7973 11253 8007
rect 11287 7973 11299 8007
rect 11241 7967 11299 7973
rect 4816 7908 5672 7936
rect 8481 7939 8539 7945
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4614 7868 4620 7880
rect 4571 7840 4620 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4816 7877 4844 7908
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 9582 7936 9588 7948
rect 8527 7908 9588 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 11256 7936 11284 7967
rect 11514 7936 11520 7948
rect 11256 7908 11520 7936
rect 11514 7896 11520 7908
rect 11572 7936 11578 7948
rect 12158 7936 12164 7948
rect 11572 7908 12164 7936
rect 11572 7896 11578 7908
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12452 7936 12480 8035
rect 12268 7908 12480 7936
rect 12621 7939 12679 7945
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5718 7868 5724 7880
rect 5031 7840 5724 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7892 7840 8033 7868
rect 7892 7828 7898 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8220 7800 8248 7831
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 8996 7840 9444 7868
rect 8996 7828 9002 7840
rect 9030 7800 9036 7812
rect 8220 7772 9036 7800
rect 9030 7760 9036 7772
rect 9088 7800 9094 7812
rect 9125 7803 9183 7809
rect 9125 7800 9137 7803
rect 9088 7772 9137 7800
rect 9088 7760 9094 7772
rect 9125 7769 9137 7772
rect 9171 7769 9183 7803
rect 9125 7763 9183 7769
rect 9306 7760 9312 7812
rect 9364 7760 9370 7812
rect 9416 7800 9444 7840
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9916 7840 10241 7868
rect 9916 7828 9922 7840
rect 10229 7837 10241 7840
rect 10275 7868 10287 7871
rect 10318 7868 10324 7880
rect 10275 7840 10324 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 10778 7868 10784 7880
rect 10459 7840 10784 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11164 7840 11713 7868
rect 9416 7772 10548 7800
rect 2590 7692 2596 7744
rect 2648 7692 2654 7744
rect 4338 7692 4344 7744
rect 4396 7692 4402 7744
rect 8386 7692 8392 7744
rect 8444 7692 8450 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 10520 7732 10548 7772
rect 10594 7760 10600 7812
rect 10652 7800 10658 7812
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 10652 7772 10701 7800
rect 10652 7760 10658 7772
rect 10689 7769 10701 7772
rect 10735 7800 10747 7803
rect 11164 7800 11192 7840
rect 11701 7837 11713 7840
rect 11747 7868 11759 7871
rect 11790 7868 11796 7880
rect 11747 7840 11796 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 12066 7868 12072 7880
rect 11931 7840 12072 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 10735 7772 11192 7800
rect 11241 7803 11299 7809
rect 10735 7769 10747 7772
rect 10689 7763 10747 7769
rect 11241 7769 11253 7803
rect 11287 7800 11299 7803
rect 11900 7800 11928 7831
rect 12066 7828 12072 7840
rect 12124 7868 12130 7880
rect 12268 7868 12296 7908
rect 12621 7905 12633 7939
rect 12667 7936 12679 7939
rect 12894 7936 12900 7948
rect 12667 7908 12900 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 12124 7840 12296 7868
rect 12124 7828 12130 7840
rect 12434 7828 12440 7880
rect 12492 7828 12498 7880
rect 11287 7772 11928 7800
rect 11287 7769 11299 7772
rect 11241 7763 11299 7769
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 12897 7803 12955 7809
rect 12897 7800 12909 7803
rect 12860 7772 12909 7800
rect 12860 7760 12866 7772
rect 12897 7769 12909 7772
rect 12943 7769 12955 7803
rect 12897 7763 12955 7769
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10520 7704 10793 7732
rect 10781 7701 10793 7704
rect 10827 7732 10839 7735
rect 11330 7732 11336 7744
rect 10827 7704 11336 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11330 7692 11336 7704
rect 11388 7732 11394 7744
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11388 7704 11805 7732
rect 11388 7692 11394 7704
rect 11793 7701 11805 7704
rect 11839 7732 11851 7735
rect 12526 7732 12532 7744
rect 11839 7704 12532 7732
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 1104 7642 14076 7664
rect 1104 7590 4918 7642
rect 4970 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 5238 7642
rect 5290 7590 10918 7642
rect 10970 7590 10982 7642
rect 11034 7590 11046 7642
rect 11098 7590 11110 7642
rect 11162 7590 11174 7642
rect 11226 7590 11238 7642
rect 11290 7590 14076 7642
rect 1104 7568 14076 7590
rect 2590 7488 2596 7540
rect 2648 7488 2654 7540
rect 3786 7488 3792 7540
rect 3844 7488 3850 7540
rect 9030 7488 9036 7540
rect 9088 7488 9094 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10284 7500 10425 7528
rect 10284 7488 10290 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11422 7528 11428 7540
rect 11112 7500 11428 7528
rect 11112 7488 11118 7500
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 12544 7500 13461 7528
rect 2308 7463 2366 7469
rect 2308 7429 2320 7463
rect 2354 7460 2366 7463
rect 2608 7460 2636 7488
rect 2354 7432 2636 7460
rect 2354 7429 2366 7432
rect 2308 7423 2366 7429
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 3804 7392 3832 7488
rect 9858 7460 9864 7472
rect 8220 7432 9864 7460
rect 3743 7364 3832 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 8220 7401 8248 7432
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8352 7364 8401 7392
rect 8352 7352 8358 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 8478 7324 8484 7336
rect 7331 7296 8484 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 2056 7188 2084 7287
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8680 7324 8708 7355
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8812 7364 8861 7392
rect 8812 7352 8818 7364
rect 8849 7361 8861 7364
rect 8895 7392 8907 7395
rect 8938 7392 8944 7404
rect 8895 7364 8944 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9508 7401 9536 7432
rect 9858 7420 9864 7432
rect 9916 7460 9922 7472
rect 9916 7432 11100 7460
rect 9916 7420 9922 7432
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9140 7324 9168 7355
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10137 7395 10195 7401
rect 10137 7392 10149 7395
rect 9732 7364 10149 7392
rect 9732 7352 9738 7364
rect 10137 7361 10149 7364
rect 10183 7361 10195 7395
rect 10594 7392 10600 7404
rect 10137 7355 10195 7361
rect 10336 7364 10600 7392
rect 8680 7296 9168 7324
rect 8772 7268 8800 7296
rect 3421 7259 3479 7265
rect 3421 7225 3433 7259
rect 3467 7256 3479 7259
rect 3878 7256 3884 7268
rect 3467 7228 3884 7256
rect 3467 7225 3479 7228
rect 3421 7219 3479 7225
rect 3878 7216 3884 7228
rect 3936 7256 3942 7268
rect 3936 7228 4752 7256
rect 3936 7216 3942 7228
rect 4724 7200 4752 7228
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7800 7228 8217 7256
rect 7800 7216 7806 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 8754 7216 8760 7268
rect 8812 7216 8818 7268
rect 9140 7256 9168 7296
rect 10336 7256 10364 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 11072 7401 11100 7432
rect 12544 7404 12572 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 12820 7432 13308 7460
rect 12820 7404 12848 7432
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 12066 7352 12072 7404
rect 12124 7352 12130 7404
rect 12526 7352 12532 7404
rect 12584 7352 12590 7404
rect 12802 7352 12808 7404
rect 12860 7352 12866 7404
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 13280 7401 13308 7432
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10468 7296 10548 7324
rect 10468 7284 10474 7296
rect 9140 7228 10364 7256
rect 10520 7256 10548 7296
rect 11330 7284 11336 7336
rect 11388 7284 11394 7336
rect 11793 7259 11851 7265
rect 11793 7256 11805 7259
rect 10520 7228 11805 7256
rect 11793 7225 11805 7228
rect 11839 7225 11851 7259
rect 11793 7219 11851 7225
rect 2406 7188 2412 7200
rect 2056 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3510 7148 3516 7200
rect 3568 7148 3574 7200
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6144 7160 6837 7188
rect 6144 7148 6150 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7190 7148 7196 7200
rect 7248 7148 7254 7200
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 7340 7160 9321 7188
rect 7340 7148 7346 7160
rect 9309 7157 9321 7160
rect 9355 7188 9367 7191
rect 9766 7188 9772 7200
rect 9355 7160 9772 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10226 7148 10232 7200
rect 10284 7148 10290 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11974 7188 11980 7200
rect 10928 7160 11980 7188
rect 10928 7148 10934 7160
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 1104 7098 14076 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 14076 7098
rect 1104 7024 14076 7046
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 4304 6956 5457 6984
rect 4304 6944 4310 6956
rect 5445 6953 5457 6956
rect 5491 6984 5503 6987
rect 5718 6984 5724 6996
rect 5491 6956 5724 6984
rect 5491 6953 5503 6956
rect 5445 6947 5503 6953
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7892 6956 8125 6984
rect 7892 6944 7898 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 8113 6947 8171 6953
rect 8128 6916 8156 6947
rect 9306 6944 9312 6996
rect 9364 6944 9370 6996
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 9493 6987 9551 6993
rect 9493 6984 9505 6987
rect 9456 6956 9505 6984
rect 9456 6944 9462 6956
rect 9493 6953 9505 6956
rect 9539 6953 9551 6987
rect 9493 6947 9551 6953
rect 10226 6944 10232 6996
rect 10284 6944 10290 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10413 6987 10471 6993
rect 10413 6984 10425 6987
rect 10376 6956 10425 6984
rect 10376 6944 10382 6956
rect 10413 6953 10425 6956
rect 10459 6953 10471 6987
rect 10413 6947 10471 6953
rect 10505 6987 10563 6993
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10870 6984 10876 6996
rect 10551 6956 10876 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11790 6984 11796 6996
rect 10980 6956 11796 6984
rect 8938 6916 8944 6928
rect 8128 6888 8944 6916
rect 8938 6876 8944 6888
rect 8996 6916 9002 6928
rect 9861 6919 9919 6925
rect 8996 6888 9812 6916
rect 8996 6876 9002 6888
rect 4062 6808 4068 6860
rect 4120 6808 4126 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 7208 6820 8493 6848
rect 7208 6792 7236 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 9232 6848 9260 6888
rect 8711 6820 9076 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 4338 6789 4344 6792
rect 4332 6780 4344 6789
rect 4299 6752 4344 6780
rect 4332 6743 4344 6752
rect 4338 6740 4344 6743
rect 4396 6740 4402 6792
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 7926 6740 7932 6792
rect 7984 6740 7990 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 5920 6644 5948 6740
rect 5997 6715 6055 6721
rect 5997 6681 6009 6715
rect 6043 6712 6055 6715
rect 6426 6715 6484 6721
rect 6426 6712 6438 6715
rect 6043 6684 6438 6712
rect 6043 6681 6055 6684
rect 5997 6675 6055 6681
rect 6426 6681 6438 6684
rect 6472 6681 6484 6715
rect 7944 6712 7972 6740
rect 6426 6675 6484 6681
rect 6564 6684 7972 6712
rect 8036 6712 8064 6743
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 8386 6712 8392 6724
rect 8036 6684 8392 6712
rect 6564 6644 6592 6684
rect 5920 6616 6592 6644
rect 7561 6647 7619 6653
rect 7561 6613 7573 6647
rect 7607 6644 7619 6647
rect 8036 6644 8064 6684
rect 8386 6672 8392 6684
rect 8444 6712 8450 6724
rect 8662 6712 8668 6724
rect 8444 6684 8668 6712
rect 8444 6672 8450 6684
rect 8662 6672 8668 6684
rect 8720 6712 8726 6724
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 8720 6684 8953 6712
rect 8720 6672 8726 6684
rect 8941 6681 8953 6684
rect 8987 6681 8999 6715
rect 9048 6712 9076 6820
rect 9140 6820 9260 6848
rect 9140 6789 9168 6820
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9498 6783 9556 6789
rect 9498 6780 9510 6783
rect 9125 6743 9183 6749
rect 9232 6752 9510 6780
rect 9232 6724 9260 6752
rect 9498 6749 9510 6752
rect 9544 6749 9556 6783
rect 9498 6743 9556 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 9214 6712 9220 6724
rect 9048 6684 9220 6712
rect 8941 6675 8999 6681
rect 7607 6616 8064 6644
rect 8956 6644 8984 6675
rect 9214 6672 9220 6684
rect 9272 6672 9278 6724
rect 9692 6712 9720 6743
rect 9784 6712 9812 6888
rect 9861 6885 9873 6919
rect 9907 6916 9919 6919
rect 10244 6916 10272 6944
rect 10594 6916 10600 6928
rect 9907 6888 10180 6916
rect 10244 6888 10600 6916
rect 9907 6885 9919 6888
rect 9861 6879 9919 6885
rect 10152 6789 10180 6888
rect 10594 6876 10600 6888
rect 10652 6916 10658 6928
rect 10781 6919 10839 6925
rect 10781 6916 10793 6919
rect 10652 6888 10793 6916
rect 10652 6876 10658 6888
rect 10781 6885 10793 6888
rect 10827 6885 10839 6919
rect 10781 6879 10839 6885
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 10686 6780 10692 6792
rect 10551 6752 10692 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 10980 6789 11008 6956
rect 11790 6944 11796 6956
rect 11848 6984 11854 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 11848 6956 13093 6984
rect 11848 6944 11854 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 11146 6916 11152 6928
rect 11072 6888 11152 6916
rect 11072 6789 11100 6888
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11422 6876 11428 6928
rect 11480 6876 11486 6928
rect 11440 6848 11468 6876
rect 11256 6820 11468 6848
rect 11256 6789 11284 6820
rect 10965 6783 11023 6789
rect 10965 6749 10977 6783
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11333 6783 11391 6789
rect 11432 6786 11490 6789
rect 11333 6749 11345 6783
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11256 6712 11284 6743
rect 9692 6684 11284 6712
rect 11348 6644 11376 6743
rect 11422 6734 11428 6786
rect 11480 6743 11490 6786
rect 11480 6734 11486 6743
rect 11974 6740 11980 6792
rect 12032 6740 12038 6792
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 11692 6715 11750 6721
rect 11692 6681 11704 6715
rect 11738 6712 11750 6715
rect 11992 6712 12020 6740
rect 11738 6684 12020 6712
rect 11738 6681 11750 6684
rect 11692 6675 11750 6681
rect 12084 6644 12112 6740
rect 8956 6616 12112 6644
rect 7607 6613 7619 6616
rect 7561 6607 7619 6613
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 1104 6554 14076 6576
rect 1104 6502 4918 6554
rect 4970 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 5238 6554
rect 5290 6502 10918 6554
rect 10970 6502 10982 6554
rect 11034 6502 11046 6554
rect 11098 6502 11110 6554
rect 11162 6502 11174 6554
rect 11226 6502 11238 6554
rect 11290 6502 14076 6554
rect 1104 6480 14076 6502
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4430 6440 4436 6452
rect 4203 6412 4436 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 7190 6440 7196 6452
rect 7024 6412 7196 6440
rect 2866 6372 2872 6384
rect 2424 6344 2872 6372
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2424 6313 2452 6344
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3044 6375 3102 6381
rect 3044 6341 3056 6375
rect 3090 6372 3102 6375
rect 3510 6372 3516 6384
rect 3090 6344 3516 6372
rect 3090 6341 3102 6344
rect 3044 6335 3102 6341
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6914 6372 6920 6384
rect 6043 6344 6920 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3602 6304 3608 6316
rect 2731 6276 3608 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 7024 6304 7052 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7282 6400 7288 6452
rect 7340 6400 7346 6452
rect 8570 6440 8576 6452
rect 8128 6412 8576 6440
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7300 6372 7328 6400
rect 7156 6344 7328 6372
rect 7377 6375 7435 6381
rect 7156 6332 7162 6344
rect 7203 6313 7231 6344
rect 7377 6341 7389 6375
rect 7423 6372 7435 6375
rect 7742 6372 7748 6384
rect 7423 6344 7748 6372
rect 7423 6341 7435 6344
rect 7377 6335 7435 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8128 6381 8156 6412
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 8754 6400 8760 6452
rect 8812 6400 8818 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 8904 6412 10916 6440
rect 8904 6400 8910 6412
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6341 8171 6375
rect 8113 6335 8171 6341
rect 8297 6375 8355 6381
rect 8297 6341 8309 6375
rect 8343 6372 8355 6375
rect 8772 6372 8800 6400
rect 8343 6344 8800 6372
rect 8343 6341 8355 6344
rect 8297 6335 8355 6341
rect 6871 6276 7052 6304
rect 7188 6307 7246 6313
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 7188 6273 7200 6307
rect 7234 6273 7246 6307
rect 7188 6267 7246 6273
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2648 6208 2789 6236
rect 2648 6196 2654 6208
rect 2777 6205 2789 6208
rect 2823 6236 2835 6239
rect 6748 6236 6776 6267
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 7006 6236 7012 6248
rect 2823 6208 2877 6236
rect 6748 6208 7012 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2792 6112 2820 6199
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7668 6236 7696 6267
rect 7116 6208 7696 6236
rect 8392 6236 8420 6267
rect 8478 6264 8484 6316
rect 8536 6307 8542 6316
rect 8573 6307 8631 6313
rect 8536 6279 8585 6307
rect 8536 6264 8542 6279
rect 8573 6273 8585 6279
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 8772 6313 8800 6344
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9674 6372 9680 6384
rect 9272 6344 9680 6372
rect 9272 6332 9278 6344
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 9950 6372 9956 6384
rect 9824 6344 9956 6372
rect 9824 6332 9830 6344
rect 9950 6332 9956 6344
rect 10008 6372 10014 6384
rect 10008 6344 10732 6372
rect 10008 6332 10014 6344
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6304 9643 6307
rect 9692 6304 9720 6332
rect 9631 6276 9720 6304
rect 9631 6273 9643 6276
rect 9585 6267 9643 6273
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10376 6276 10425 6304
rect 10376 6264 10382 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10704 6313 10732 6344
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 8392 6208 9076 6236
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 4120 6140 4752 6168
rect 4120 6128 4126 6140
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1820 6072 2053 6100
rect 1820 6060 1826 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 4080 6100 4108 6128
rect 4724 6109 4752 6140
rect 6638 6128 6644 6180
rect 6696 6168 6702 6180
rect 7116 6168 7144 6208
rect 6696 6140 7144 6168
rect 6696 6128 6702 6140
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 7929 6171 7987 6177
rect 7929 6168 7941 6171
rect 7800 6140 7941 6168
rect 7800 6128 7806 6140
rect 7929 6137 7941 6140
rect 7975 6168 7987 6171
rect 8386 6168 8392 6180
rect 7975 6140 8392 6168
rect 7975 6137 7987 6140
rect 7929 6131 7987 6137
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 9048 6168 9076 6208
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10134 6236 10140 6248
rect 9548 6208 10140 6236
rect 9548 6196 9554 6208
rect 10134 6196 10140 6208
rect 10192 6236 10198 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10192 6208 10793 6236
rect 10192 6196 10198 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 10888 6236 10916 6412
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11388 6412 11897 6440
rect 11388 6400 11394 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 11532 6344 12112 6372
rect 11532 6316 11560 6344
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 11112 6276 11161 6304
rect 11112 6264 11118 6276
rect 11149 6273 11161 6276
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 11514 6264 11520 6316
rect 11572 6264 11578 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 12084 6313 12112 6344
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12894 6304 12900 6316
rect 12575 6276 12900 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 11900 6236 11928 6264
rect 10888 6208 11928 6236
rect 12253 6239 12311 6245
rect 10042 6168 10048 6180
rect 9048 6140 10048 6168
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 2832 6072 4108 6100
rect 4709 6103 4767 6109
rect 2832 6060 2838 6072
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 6178 6100 6184 6112
rect 4755 6072 6184 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7006 6060 7012 6112
rect 7064 6060 7070 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8846 6100 8852 6112
rect 7616 6072 8852 6100
rect 7616 6060 7622 6072
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 9122 6060 9128 6112
rect 9180 6060 9186 6112
rect 9214 6060 9220 6112
rect 9272 6060 9278 6112
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 10888 6109 10916 6208
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12802 6236 12808 6248
rect 12299 6208 12808 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 11057 6171 11115 6177
rect 11057 6137 11069 6171
rect 11103 6168 11115 6171
rect 11422 6168 11428 6180
rect 11103 6140 11428 6168
rect 11103 6137 11115 6140
rect 11057 6131 11115 6137
rect 11422 6128 11428 6140
rect 11480 6128 11486 6180
rect 10873 6103 10931 6109
rect 10873 6069 10885 6103
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 11241 6103 11299 6109
rect 11241 6069 11253 6103
rect 11287 6100 11299 6103
rect 11330 6100 11336 6112
rect 11287 6072 11336 6100
rect 11287 6069 11299 6072
rect 11241 6063 11299 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12066 6060 12072 6112
rect 12124 6060 12130 6112
rect 1104 6010 14076 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 14076 6010
rect 1104 5936 14076 5958
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 2556 5868 3065 5896
rect 2556 5856 2562 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 6178 5896 6184 5908
rect 3053 5859 3111 5865
rect 5460 5868 6184 5896
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4212 5800 5120 5828
rect 4212 5788 4218 5800
rect 3528 5732 4108 5760
rect 3528 5701 3556 5732
rect 4080 5704 4108 5732
rect 4356 5732 5028 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1848 5695 1906 5701
rect 1848 5661 1860 5695
rect 1894 5661 1906 5695
rect 1848 5655 1906 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 1596 5556 1624 5655
rect 1762 5584 1768 5636
rect 1820 5624 1826 5636
rect 1872 5624 1900 5655
rect 1820 5596 1900 5624
rect 3252 5624 3280 5655
rect 3988 5624 4016 5655
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4120 5664 4261 5692
rect 4120 5652 4126 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4356 5636 4384 5732
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4798 5692 4804 5704
rect 4755 5664 4804 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5000 5701 5028 5732
rect 5092 5701 5120 5800
rect 5460 5769 5488 5868
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 7006 5856 7012 5908
rect 7064 5856 7070 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8036 5868 9137 5896
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 7024 5692 7052 5856
rect 5077 5655 5135 5661
rect 5184 5664 7052 5692
rect 7101 5695 7159 5701
rect 3252 5596 4292 5624
rect 1820 5584 1826 5596
rect 2774 5556 2780 5568
rect 1596 5528 2780 5556
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3016 5528 3433 5556
rect 3016 5516 3022 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 3421 5519 3479 5525
rect 3786 5516 3792 5568
rect 3844 5516 3850 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4264 5556 4292 5596
rect 4338 5584 4344 5636
rect 4396 5584 4402 5636
rect 4908 5624 4936 5655
rect 5184 5624 5212 5664
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7190 5692 7196 5704
rect 7147 5664 7196 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7742 5692 7748 5704
rect 7331 5664 7748 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 4908 5596 5212 5624
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5690 5627 5748 5633
rect 5690 5624 5702 5627
rect 5399 5596 5702 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5690 5593 5702 5596
rect 5736 5593 5748 5627
rect 5690 5587 5748 5593
rect 6638 5584 6644 5636
rect 6696 5584 6702 5636
rect 7208 5624 7236 5652
rect 8036 5624 8064 5868
rect 9125 5865 9137 5868
rect 9171 5896 9183 5899
rect 9490 5896 9496 5908
rect 9171 5868 9496 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10318 5896 10324 5908
rect 9916 5868 10324 5896
rect 9916 5856 9922 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 8570 5788 8576 5840
rect 8628 5788 8634 5840
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 8812 5800 9260 5828
rect 8812 5788 8818 5800
rect 8588 5692 8616 5788
rect 9232 5769 9260 5800
rect 9398 5788 9404 5840
rect 9456 5828 9462 5840
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 9456 5800 10057 5828
rect 9456 5788 9462 5800
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10045 5791 10103 5797
rect 10137 5831 10195 5837
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10594 5828 10600 5840
rect 10183 5800 10600 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10594 5788 10600 5800
rect 10652 5828 10658 5840
rect 11698 5828 11704 5840
rect 10652 5800 11704 5828
rect 10652 5788 10658 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5760 9275 5763
rect 9263 5732 9674 5760
rect 9263 5729 9275 5732
rect 9217 5723 9275 5729
rect 9030 5692 9036 5704
rect 8588 5664 9036 5692
rect 9030 5652 9036 5664
rect 9088 5692 9094 5704
rect 9493 5695 9551 5701
rect 9493 5692 9505 5695
rect 9088 5664 9505 5692
rect 9088 5652 9094 5664
rect 9493 5661 9505 5664
rect 9539 5661 9551 5695
rect 9646 5692 9674 5732
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9646 5664 9965 5692
rect 9493 5655 9551 5661
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10376 5664 10425 5692
rect 10376 5652 10382 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 6840 5596 7144 5624
rect 7208 5596 8064 5624
rect 8128 5596 9904 5624
rect 6656 5556 6684 5584
rect 6840 5565 6868 5596
rect 4264 5528 6684 5556
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5525 6883 5559
rect 6825 5519 6883 5525
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 7116 5556 7144 5596
rect 7374 5556 7380 5568
rect 7116 5528 7380 5556
rect 7374 5516 7380 5528
rect 7432 5556 7438 5568
rect 8128 5556 8156 5596
rect 9876 5568 9904 5596
rect 7432 5528 8156 5556
rect 7432 5516 7438 5528
rect 8938 5516 8944 5568
rect 8996 5516 9002 5568
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 9858 5516 9864 5568
rect 9916 5516 9922 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11514 5556 11520 5568
rect 11296 5528 11520 5556
rect 11296 5516 11302 5528
rect 11514 5516 11520 5528
rect 11572 5556 11578 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11572 5528 11805 5556
rect 11572 5516 11578 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 1104 5466 14076 5488
rect 1104 5414 4918 5466
rect 4970 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 5238 5466
rect 5290 5414 10918 5466
rect 10970 5414 10982 5466
rect 11034 5414 11046 5466
rect 11098 5414 11110 5466
rect 11162 5414 11174 5466
rect 11226 5414 11238 5466
rect 11290 5414 14076 5466
rect 1104 5392 14076 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 2924 5324 3372 5352
rect 2924 5312 2930 5324
rect 2624 5287 2682 5293
rect 2624 5253 2636 5287
rect 2670 5284 2682 5287
rect 2961 5287 3019 5293
rect 2961 5284 2973 5287
rect 2670 5256 2973 5284
rect 2670 5253 2682 5256
rect 2624 5247 2682 5253
rect 2961 5253 2973 5256
rect 3007 5253 3019 5287
rect 2961 5247 3019 5253
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2832 5188 2881 5216
rect 2832 5176 2838 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3234 5176 3240 5228
rect 3292 5176 3298 5228
rect 3344 5225 3372 5324
rect 3786 5312 3792 5364
rect 3844 5312 3850 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 7098 5352 7104 5364
rect 4120 5324 7104 5352
rect 4120 5312 4126 5324
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 9122 5312 9128 5364
rect 9180 5312 9186 5364
rect 9762 5355 9820 5361
rect 9762 5321 9774 5355
rect 9808 5352 9820 5355
rect 9808 5324 10180 5352
rect 9808 5321 9820 5324
rect 9762 5315 9820 5321
rect 3804 5284 3832 5312
rect 9140 5284 9168 5312
rect 10152 5284 10180 5324
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10284 5324 10425 5352
rect 10284 5312 10290 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10520 5324 11560 5352
rect 10520 5284 10548 5324
rect 11532 5284 11560 5324
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 11762 5287 11820 5293
rect 11762 5284 11774 5287
rect 3436 5256 3832 5284
rect 3896 5256 4660 5284
rect 9140 5256 9628 5284
rect 3436 5225 3464 5256
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3344 5148 3372 5179
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3786 5216 3792 5228
rect 3660 5188 3792 5216
rect 3660 5176 3666 5188
rect 3786 5176 3792 5188
rect 3844 5216 3850 5228
rect 3896 5216 3924 5256
rect 3844 5188 3924 5216
rect 3844 5176 3850 5188
rect 4246 5176 4252 5228
rect 4304 5176 4310 5228
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 4632 5225 4660 5256
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 4798 5216 4804 5228
rect 4663 5188 4804 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4798 5176 4804 5188
rect 4856 5216 4862 5228
rect 5442 5216 5448 5228
rect 4856 5188 5448 5216
rect 4856 5176 4862 5188
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 6914 5216 6920 5228
rect 6687 5188 6920 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9088 5188 9321 5216
rect 9088 5176 9094 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9600 5225 9628 5256
rect 9692 5256 9996 5284
rect 10152 5256 10548 5284
rect 10612 5256 11468 5284
rect 11532 5256 11774 5284
rect 9692 5228 9720 5256
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 9456 5188 9505 5216
rect 9456 5176 9462 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 4062 5148 4068 5160
rect 3344 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5148 4126 5160
rect 4356 5148 4384 5176
rect 4120 5120 4384 5148
rect 4120 5108 4126 5120
rect 9600 5080 9628 5179
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 9968 5225 9996 5256
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 9876 5148 9904 5179
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 10612 5225 10640 5256
rect 11440 5228 11468 5256
rect 11762 5253 11774 5256
rect 11808 5253 11820 5287
rect 11762 5247 11820 5253
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11330 5216 11336 5228
rect 10827 5188 11336 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11422 5176 11428 5228
rect 11480 5176 11486 5228
rect 10229 5151 10287 5157
rect 9876 5120 10180 5148
rect 10152 5089 10180 5120
rect 10229 5117 10241 5151
rect 10275 5148 10287 5151
rect 10336 5148 10364 5176
rect 10275 5120 10364 5148
rect 10428 5148 10456 5176
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10428 5120 10701 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 10919 5120 11376 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 3436 5052 4200 5080
rect 9600 5052 10057 5080
rect 1489 5015 1547 5021
rect 1489 4981 1501 5015
rect 1535 5012 1547 5015
rect 1578 5012 1584 5024
rect 1535 4984 1584 5012
rect 1535 4981 1547 4984
rect 1489 4975 1547 4981
rect 1578 4972 1584 4984
rect 1636 5012 1642 5024
rect 3436 5012 3464 5052
rect 4172 5024 4200 5052
rect 10045 5049 10057 5052
rect 10091 5049 10103 5083
rect 10045 5043 10103 5049
rect 10137 5083 10195 5089
rect 10137 5049 10149 5083
rect 10183 5049 10195 5083
rect 10137 5043 10195 5049
rect 11348 5024 11376 5120
rect 11514 5108 11520 5160
rect 11572 5108 11578 5160
rect 1636 4984 3464 5012
rect 1636 4972 1642 4984
rect 3970 4972 3976 5024
rect 4028 4972 4034 5024
rect 4154 4972 4160 5024
rect 4212 4972 4218 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 5592 4984 6469 5012
rect 5592 4972 5598 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 9493 5015 9551 5021
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 10226 5012 10232 5024
rect 9539 4984 10232 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 11330 4972 11336 5024
rect 11388 4972 11394 5024
rect 1104 4922 14076 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 14076 4922
rect 1104 4848 14076 4870
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 8938 4808 8944 4820
rect 8628 4780 8944 4808
rect 8628 4768 8634 4780
rect 8938 4768 8944 4780
rect 8996 4808 9002 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8996 4780 9321 4808
rect 8996 4768 9002 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9309 4771 9367 4777
rect 9674 4768 9680 4820
rect 9732 4768 9738 4820
rect 10410 4808 10416 4820
rect 9784 4780 10416 4808
rect 4080 4672 4108 4768
rect 5534 4672 5540 4684
rect 4080 4644 5540 4672
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4356 4613 4384 4644
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3844 4576 4077 4604
rect 3844 4564 3850 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4522 4604 4528 4616
rect 4479 4576 4528 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4264 4536 4292 4567
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 5184 4613 5212 4644
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4764 4576 5089 4604
rect 4764 4564 4770 4576
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 4614 4536 4620 4548
rect 4264 4508 4620 4536
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 5276 4536 5304 4567
rect 5442 4564 5448 4616
rect 5500 4564 5506 4616
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 8904 4576 9229 4604
rect 8904 4564 8910 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 9784 4604 9812 4780
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10226 4700 10232 4752
rect 10284 4700 10290 4752
rect 9539 4576 9812 4604
rect 9861 4607 9919 4613
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 6362 4536 6368 4548
rect 5276 4508 6368 4536
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 9876 4536 9904 4567
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 10008 4576 10057 4604
rect 10008 4564 10014 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10134 4564 10140 4616
rect 10192 4564 10198 4616
rect 10244 4613 10272 4700
rect 10318 4632 10324 4684
rect 10376 4632 10382 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 11572 4644 11928 4672
rect 11572 4632 11578 4644
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10336 4536 10364 4632
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 11790 4604 11796 4616
rect 10459 4576 11796 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 11900 4604 11928 4644
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 11900 4576 13553 4604
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13296 4539 13354 4545
rect 9732 4508 10364 4536
rect 10428 4508 12204 4536
rect 9732 4496 9738 4508
rect 4706 4428 4712 4480
rect 4764 4428 4770 4480
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 9214 4468 9220 4480
rect 8444 4440 9220 4468
rect 8444 4428 8450 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 10428 4468 10456 4508
rect 9640 4440 10456 4468
rect 10597 4471 10655 4477
rect 9640 4428 9646 4440
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 10686 4468 10692 4480
rect 10643 4440 10692 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 12176 4477 12204 4508
rect 13296 4505 13308 4539
rect 13342 4536 13354 4539
rect 13446 4536 13452 4548
rect 13342 4508 13452 4536
rect 13342 4505 13354 4508
rect 13296 4499 13354 4505
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4437 12219 4471
rect 12161 4431 12219 4437
rect 1104 4378 14076 4400
rect 1104 4326 4918 4378
rect 4970 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 5238 4378
rect 5290 4326 10918 4378
rect 10970 4326 10982 4378
rect 11034 4326 11046 4378
rect 11098 4326 11110 4378
rect 11162 4326 11174 4378
rect 11226 4326 11238 4378
rect 11290 4326 14076 4378
rect 1104 4304 14076 4326
rect 2866 4224 2872 4276
rect 2924 4224 2930 4276
rect 3694 4224 3700 4276
rect 3752 4224 3758 4276
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 6362 4224 6368 4276
rect 6420 4224 6426 4276
rect 7098 4224 7104 4276
rect 7156 4224 7162 4276
rect 8570 4264 8576 4276
rect 8220 4236 8576 4264
rect 2884 4196 2912 4224
rect 2884 4168 3188 4196
rect 2774 4088 2780 4140
rect 2832 4088 2838 4140
rect 3050 4088 3056 4140
rect 3108 4088 3114 4140
rect 3160 4137 3188 4168
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3712 4128 3740 4224
rect 3780 4199 3838 4205
rect 3780 4165 3792 4199
rect 3826 4196 3838 4199
rect 3970 4196 3976 4208
rect 3826 4168 3976 4196
rect 3826 4165 3838 4168
rect 3780 4159 3838 4165
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 5552 4196 5580 4224
rect 5552 4168 5764 4196
rect 3467 4100 3740 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5500 4100 5580 4128
rect 5500 4088 5506 4100
rect 2792 4060 2820 4088
rect 3510 4060 3516 4072
rect 2792 4032 3516 4060
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 5552 3992 5580 4100
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 5736 4137 5764 4168
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6638 4128 6644 4140
rect 6595 4100 6644 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6748 4060 6776 4091
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7116 4128 7144 4224
rect 8220 4205 8248 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 9674 4264 9680 4276
rect 8680 4236 9680 4264
rect 7561 4199 7619 4205
rect 7561 4165 7573 4199
rect 7607 4196 7619 4199
rect 8205 4199 8263 4205
rect 7607 4168 8156 4196
rect 7607 4165 7619 4168
rect 7561 4159 7619 4165
rect 6880 4100 7144 4128
rect 6880 4088 6886 4100
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8128 4128 8156 4168
rect 8205 4165 8217 4199
rect 8251 4165 8263 4199
rect 8680 4196 8708 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 13446 4224 13452 4276
rect 13504 4264 13510 4276
rect 13541 4267 13599 4273
rect 13541 4264 13553 4267
rect 13504 4236 13553 4264
rect 13504 4224 13510 4236
rect 13541 4233 13553 4236
rect 13587 4233 13599 4267
rect 13541 4227 13599 4233
rect 8205 4159 8263 4165
rect 8312 4168 8708 4196
rect 8312 4137 8340 4168
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 11514 4196 11520 4208
rect 10008 4168 11520 4196
rect 10008 4156 10014 4168
rect 11514 4156 11520 4168
rect 11572 4196 11578 4208
rect 11572 4168 12204 4196
rect 11572 4156 11578 4168
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8128 4100 8309 4128
rect 8021 4091 8079 4097
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 7300 4060 7328 4088
rect 8036 4060 8064 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8711 4100 8800 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 6748 4032 7328 4060
rect 7852 4032 8064 4060
rect 8404 4060 8432 4088
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8404 4032 8585 4060
rect 5552 3964 7512 3992
rect 7484 3936 7512 3964
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 2648 3896 2789 3924
rect 2648 3884 2654 3896
rect 2777 3893 2789 3896
rect 2823 3893 2835 3927
rect 2777 3887 2835 3893
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4304 3896 4905 3924
rect 4304 3884 4310 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 4893 3887 4951 3893
rect 6089 3927 6147 3933
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 6178 3924 6184 3936
rect 6135 3896 6184 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 7466 3884 7472 3936
rect 7524 3884 7530 3936
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 7852 3924 7880 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 8772 4060 8800 4100
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8996 4100 9137 4128
rect 8996 4088 9002 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 12176 4137 12204 4168
rect 10209 4131 10267 4137
rect 10209 4128 10221 4131
rect 9824 4100 10221 4128
rect 9824 4088 9830 4100
rect 10209 4097 10221 4100
rect 10255 4097 10267 4131
rect 10209 4091 10267 4097
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12428 4131 12486 4137
rect 12428 4097 12440 4131
rect 12474 4128 12486 4131
rect 13538 4128 13544 4140
rect 12474 4100 13544 4128
rect 12474 4097 12486 4100
rect 12428 4091 12486 4097
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 8772 4032 9352 4060
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8772 3992 8800 4032
rect 9324 4001 9352 4032
rect 9950 4020 9956 4072
rect 10008 4020 10014 4072
rect 7975 3964 8800 3992
rect 9309 3995 9367 4001
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 8938 3924 8944 3936
rect 7852 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9030 3884 9036 3936
rect 9088 3884 9094 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12066 3924 12072 3936
rect 11388 3896 12072 3924
rect 11388 3884 11394 3896
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 1104 3834 14076 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 14076 3834
rect 1104 3760 14076 3782
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4430 3720 4436 3732
rect 4387 3692 4436 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 5859 3692 7328 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 7300 3664 7328 3692
rect 11790 3680 11796 3732
rect 11848 3720 11854 3732
rect 12158 3720 12164 3732
rect 11848 3692 12164 3720
rect 11848 3680 11854 3692
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 7282 3612 7288 3664
rect 7340 3612 7346 3664
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 4062 3584 4068 3596
rect 3568 3556 4068 3584
rect 3568 3544 3574 3556
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4120 3556 4445 3584
rect 4120 3544 4126 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 3528 3516 3556 3544
rect 2271 3488 3556 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 3878 3476 3884 3528
rect 3936 3476 3942 3528
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 4448 3516 4476 3547
rect 6178 3525 6184 3528
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 4448 3488 5917 3516
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 6172 3516 6184 3525
rect 6139 3488 6184 3516
rect 5905 3479 5963 3485
rect 6172 3479 6184 3488
rect 6178 3476 6184 3479
rect 6236 3476 6242 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 7423 3488 8953 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 8941 3485 8953 3488
rect 8987 3516 8999 3519
rect 9950 3516 9956 3528
rect 8987 3488 9956 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9950 3476 9956 3488
rect 10008 3516 10014 3528
rect 10686 3525 10692 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10008 3488 10425 3516
rect 10008 3476 10014 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10680 3516 10692 3525
rect 10647 3488 10692 3516
rect 10413 3479 10471 3485
rect 10680 3479 10692 3488
rect 10686 3476 10692 3479
rect 10744 3476 10750 3528
rect 2492 3451 2550 3457
rect 2492 3417 2504 3451
rect 2538 3448 2550 3451
rect 2590 3448 2596 3460
rect 2538 3420 2596 3448
rect 2538 3417 2550 3420
rect 2492 3411 2550 3417
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 3973 3451 4031 3457
rect 3973 3417 3985 3451
rect 4019 3448 4031 3451
rect 4264 3448 4292 3476
rect 4019 3420 4292 3448
rect 4700 3451 4758 3457
rect 4019 3417 4031 3420
rect 3973 3411 4031 3417
rect 4700 3417 4712 3451
rect 4746 3448 4758 3451
rect 4798 3448 4804 3460
rect 4746 3420 4804 3448
rect 4746 3417 4758 3420
rect 4700 3411 4758 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 7644 3451 7702 3457
rect 7644 3417 7656 3451
rect 7690 3448 7702 3451
rect 7742 3448 7748 3460
rect 7690 3420 7748 3448
rect 7690 3417 7702 3420
rect 7644 3411 7702 3417
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8846 3448 8852 3460
rect 8720 3420 8852 3448
rect 8720 3408 8726 3420
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9186 3451 9244 3457
rect 9186 3448 9198 3451
rect 9088 3420 9198 3448
rect 9088 3408 9094 3420
rect 9186 3417 9198 3420
rect 9232 3417 9244 3451
rect 9186 3411 9244 3417
rect 3602 3340 3608 3392
rect 3660 3340 3666 3392
rect 7285 3383 7343 3389
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7558 3380 7564 3392
rect 7331 3352 7564 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 8864 3380 8892 3408
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 8864 3352 10333 3380
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 10321 3343 10379 3349
rect 1104 3290 14076 3312
rect 1104 3238 4918 3290
rect 4970 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 5238 3290
rect 5290 3238 10918 3290
rect 10970 3238 10982 3290
rect 11034 3238 11046 3290
rect 11098 3238 11110 3290
rect 11162 3238 11174 3290
rect 11226 3238 11238 3290
rect 11290 3238 14076 3290
rect 1104 3216 14076 3238
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3234 3176 3240 3188
rect 3099 3148 3240 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3602 3176 3608 3188
rect 3467 3148 3608 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5684 3148 6377 3176
rect 5684 3136 5690 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 7558 3176 7564 3188
rect 6779 3148 7564 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 8662 3136 8668 3188
rect 8720 3136 8726 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 8938 3136 8944 3188
rect 8996 3136 9002 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 4154 3108 4160 3120
rect 3252 3080 4160 3108
rect 3252 3049 3280 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 4862 3111 4920 3117
rect 4862 3108 4874 3111
rect 4764 3080 4874 3108
rect 4764 3068 4770 3080
rect 4862 3077 4874 3080
rect 4908 3077 4920 3111
rect 4862 3071 4920 3077
rect 6822 3068 6828 3120
rect 6880 3068 6886 3120
rect 8481 3111 8539 3117
rect 8481 3077 8493 3111
rect 8527 3108 8539 3111
rect 8570 3108 8576 3120
rect 8527 3080 8576 3108
rect 8527 3077 8539 3080
rect 8481 3071 8539 3077
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 6822 3065 6880 3068
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3878 3040 3884 3052
rect 3559 3012 3884 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4120 3012 4629 3040
rect 4120 3000 4126 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6638 3040 6644 3052
rect 6595 3012 6644 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6822 3031 6834 3065
rect 6868 3031 6880 3065
rect 8772 3049 8800 3136
rect 6822 3025 6880 3031
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3040 8815 3043
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8803 3012 8861 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9999 3012 10241 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10229 3009 10241 3012
rect 10275 3040 10287 3043
rect 10336 3040 10364 3136
rect 10275 3012 10364 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 8478 2864 8484 2916
rect 8536 2864 8542 2916
rect 5994 2796 6000 2848
rect 6052 2796 6058 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 1104 2746 14076 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 14076 2746
rect 1104 2672 14076 2694
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4672 2604 4997 2632
rect 4672 2592 4678 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 6638 2592 6644 2644
rect 6696 2592 6702 2644
rect 13538 2592 13544 2644
rect 13596 2592 13602 2644
rect 4154 2524 4160 2576
rect 4212 2564 4218 2576
rect 6656 2564 6684 2592
rect 4212 2536 6684 2564
rect 4212 2524 4218 2536
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 2958 2428 2964 2440
rect 2547 2400 2964 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3476 2400 3985 2428
rect 3476 2388 3482 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 5184 2437 5212 2536
rect 5994 2496 6000 2508
rect 5368 2468 6000 2496
rect 5368 2437 5396 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4304 2400 4905 2428
rect 4304 2388 4310 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2397 5503 2431
rect 6012 2428 6040 2456
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 6012 2400 6101 2428
rect 5445 2391 5503 2397
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 5460 2360 5488 2391
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 7282 2388 7288 2440
rect 7340 2388 7346 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 7616 2400 8493 2428
rect 7616 2388 7622 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9858 2428 9864 2440
rect 9723 2400 9864 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10468 2400 10885 2428
rect 10468 2388 10474 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12216 2400 13277 2428
rect 12216 2388 12222 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 14182 2428 14188 2440
rect 13771 2400 14188 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 6840 2360 6868 2388
rect 5460 2332 6868 2360
rect 1026 2252 1032 2304
rect 1084 2292 1090 2304
rect 1397 2295 1455 2301
rect 1397 2292 1409 2295
rect 1084 2264 1409 2292
rect 1084 2252 1090 2264
rect 1397 2261 1409 2264
rect 1443 2261 1455 2295
rect 1397 2255 1455 2261
rect 2314 2252 2320 2304
rect 2372 2252 2378 2304
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3476 2264 3801 2292
rect 3476 2252 3482 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 4706 2252 4712 2304
rect 4764 2252 4770 2304
rect 5902 2252 5908 2304
rect 5960 2252 5966 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8260 2264 8309 2292
rect 8260 2252 8266 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 9490 2252 9496 2304
rect 9548 2252 9554 2304
rect 10686 2252 10692 2304
rect 10744 2252 10750 2304
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 1104 2202 14076 2224
rect 1104 2150 4918 2202
rect 4970 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 5238 2202
rect 5290 2150 10918 2202
rect 10970 2150 10982 2202
rect 11034 2150 11046 2202
rect 11098 2150 11110 2202
rect 11162 2150 11174 2202
rect 11226 2150 11238 2202
rect 11290 2150 14076 2202
rect 1104 2128 14076 2150
<< via1 >>
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 1032 14560 1084 14612
rect 2320 14560 2372 14612
rect 3056 14560 3108 14612
rect 4068 14560 4120 14612
rect 5080 14560 5132 14612
rect 6092 14560 6144 14612
rect 7104 14560 7156 14612
rect 7840 14560 7892 14612
rect 9128 14560 9180 14612
rect 2504 14356 2556 14408
rect 3516 14356 3568 14408
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4436 14356 4488 14408
rect 5724 14356 5776 14408
rect 6920 14356 6972 14408
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 9404 14399 9456 14408
rect 9404 14365 9413 14399
rect 9413 14365 9447 14399
rect 9447 14365 9456 14399
rect 9404 14356 9456 14365
rect 11152 14356 11204 14408
rect 12164 14356 12216 14408
rect 13176 14356 13228 14408
rect 5448 14288 5500 14340
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 13268 14220 13320 14272
rect 4918 14118 4970 14170
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 5238 14118 5290 14170
rect 10918 14118 10970 14170
rect 10982 14118 11034 14170
rect 11046 14118 11098 14170
rect 11110 14118 11162 14170
rect 11174 14118 11226 14170
rect 11238 14118 11290 14170
rect 5356 13880 5408 13932
rect 5448 13880 5500 13932
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 9772 13880 9824 13932
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 4528 13744 4580 13796
rect 5264 13744 5316 13796
rect 10692 13744 10744 13796
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 4160 13676 4212 13728
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 6368 13676 6420 13685
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 9404 13676 9456 13728
rect 11336 13676 11388 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 5264 13472 5316 13524
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 4988 13404 5040 13456
rect 8392 13472 8444 13524
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 9680 13472 9732 13524
rect 9956 13472 10008 13524
rect 2136 13268 2188 13320
rect 2872 13268 2924 13320
rect 2320 13243 2372 13252
rect 2320 13209 2354 13243
rect 2354 13209 2372 13243
rect 2320 13200 2372 13209
rect 4160 13200 4212 13252
rect 9680 13268 9732 13320
rect 10324 13268 10376 13320
rect 6368 13200 6420 13252
rect 7656 13200 7708 13252
rect 8300 13200 8352 13252
rect 10232 13200 10284 13252
rect 5448 13132 5500 13184
rect 6920 13132 6972 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 10692 13132 10744 13184
rect 11612 13132 11664 13184
rect 12072 13132 12124 13184
rect 12256 13200 12308 13252
rect 12348 13132 12400 13184
rect 4918 13030 4970 13082
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 5238 13030 5290 13082
rect 10918 13030 10970 13082
rect 10982 13030 11034 13082
rect 11046 13030 11098 13082
rect 11110 13030 11162 13082
rect 11174 13030 11226 13082
rect 11238 13030 11290 13082
rect 2320 12928 2372 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 7104 12928 7156 12980
rect 7196 12928 7248 12980
rect 7656 12971 7708 12980
rect 7656 12937 7665 12971
rect 7665 12937 7699 12971
rect 7699 12937 7708 12971
rect 7656 12928 7708 12937
rect 9680 12928 9732 12980
rect 2136 12860 2188 12912
rect 2228 12792 2280 12844
rect 4896 12860 4948 12912
rect 2964 12792 3016 12844
rect 4068 12724 4120 12776
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 4620 12656 4672 12708
rect 5172 12724 5224 12776
rect 3332 12588 3384 12640
rect 3792 12588 3844 12640
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 6920 12792 6972 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7012 12656 7064 12708
rect 6828 12588 6880 12640
rect 7656 12588 7708 12640
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 9220 12860 9272 12912
rect 9312 12860 9364 12912
rect 9864 12860 9916 12912
rect 9956 12860 10008 12912
rect 11244 12928 11296 12980
rect 10600 12792 10652 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 10784 12792 10836 12844
rect 11336 12860 11388 12912
rect 9312 12724 9364 12776
rect 9128 12656 9180 12708
rect 10508 12724 10560 12776
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 12072 12928 12124 12980
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12348 12792 12400 12844
rect 11612 12724 11664 12776
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 12716 12724 12768 12776
rect 12164 12656 12216 12708
rect 8484 12588 8536 12640
rect 9680 12588 9732 12640
rect 10784 12588 10836 12640
rect 11244 12588 11296 12640
rect 11336 12588 11388 12640
rect 12256 12588 12308 12640
rect 12532 12588 12584 12640
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 2320 12384 2372 12436
rect 3700 12384 3752 12436
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 5172 12384 5224 12436
rect 3424 12316 3476 12368
rect 2964 12155 3016 12164
rect 2964 12121 2973 12155
rect 2973 12121 3007 12155
rect 3007 12121 3016 12155
rect 2964 12112 3016 12121
rect 4896 12316 4948 12368
rect 5356 12316 5408 12368
rect 3792 12248 3844 12300
rect 5448 12248 5500 12300
rect 5540 12248 5592 12300
rect 3608 12180 3660 12232
rect 3884 12180 3936 12232
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 4252 12180 4304 12232
rect 4528 12180 4580 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 5540 12112 5592 12164
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 6552 12384 6604 12436
rect 6736 12384 6788 12436
rect 8392 12384 8444 12436
rect 10324 12384 10376 12436
rect 10416 12384 10468 12436
rect 6920 12316 6972 12368
rect 10784 12316 10836 12368
rect 11612 12384 11664 12436
rect 11704 12384 11756 12436
rect 11244 12316 11296 12368
rect 7012 12180 7064 12232
rect 10140 12248 10192 12300
rect 11520 12316 11572 12368
rect 11888 12359 11940 12368
rect 11888 12325 11897 12359
rect 11897 12325 11931 12359
rect 11931 12325 11940 12359
rect 11888 12316 11940 12325
rect 11980 12316 12032 12368
rect 7564 12180 7616 12232
rect 3700 12044 3752 12096
rect 4620 12044 4672 12096
rect 4896 12044 4948 12096
rect 7288 12112 7340 12164
rect 8484 12180 8536 12232
rect 9128 12180 9180 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10232 12180 10284 12232
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 10876 12180 10928 12232
rect 11152 12180 11204 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 11888 12180 11940 12232
rect 11428 12155 11480 12164
rect 11428 12121 11437 12155
rect 11437 12121 11471 12155
rect 11471 12121 11480 12155
rect 11428 12112 11480 12121
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 12440 12180 12492 12232
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 7012 12044 7064 12096
rect 8116 12044 8168 12096
rect 9864 12044 9916 12096
rect 10508 12044 10560 12096
rect 10876 12044 10928 12096
rect 12256 12044 12308 12096
rect 12440 12087 12492 12096
rect 12440 12053 12455 12087
rect 12455 12053 12489 12087
rect 12489 12053 12492 12087
rect 12440 12044 12492 12053
rect 12716 12112 12768 12164
rect 12808 12044 12860 12096
rect 4918 11942 4970 11994
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 5238 11942 5290 11994
rect 10918 11942 10970 11994
rect 10982 11942 11034 11994
rect 11046 11942 11098 11994
rect 11110 11942 11162 11994
rect 11174 11942 11226 11994
rect 11238 11942 11290 11994
rect 2964 11840 3016 11892
rect 3608 11840 3660 11892
rect 4528 11883 4580 11892
rect 4528 11849 4537 11883
rect 4537 11849 4571 11883
rect 4571 11849 4580 11883
rect 4528 11840 4580 11849
rect 7564 11840 7616 11892
rect 7656 11840 7708 11892
rect 4068 11704 4120 11756
rect 4620 11704 4672 11756
rect 4896 11704 4948 11756
rect 5816 11772 5868 11824
rect 6368 11704 6420 11756
rect 7012 11704 7064 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7932 11840 7984 11892
rect 9772 11840 9824 11892
rect 10048 11840 10100 11892
rect 9864 11772 9916 11824
rect 3056 11636 3108 11688
rect 2964 11500 3016 11552
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 3884 11636 3936 11688
rect 7104 11636 7156 11688
rect 9772 11704 9824 11756
rect 11520 11840 11572 11892
rect 11612 11840 11664 11892
rect 12348 11840 12400 11892
rect 12440 11840 12492 11892
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 10140 11704 10192 11756
rect 10692 11704 10744 11756
rect 11980 11704 12032 11756
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 10416 11636 10468 11688
rect 10508 11636 10560 11688
rect 10784 11636 10836 11688
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 4712 11500 4764 11552
rect 7380 11500 7432 11552
rect 10600 11568 10652 11620
rect 11336 11500 11388 11552
rect 11704 11500 11756 11552
rect 13176 11500 13228 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 2504 11296 2556 11348
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 3332 11092 3384 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4252 11296 4304 11348
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 3700 11160 3752 11212
rect 5356 11228 5408 11280
rect 7932 11228 7984 11280
rect 11796 11296 11848 11348
rect 12440 11296 12492 11348
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 4252 11092 4304 11144
rect 9404 11160 9456 11212
rect 10232 11228 10284 11280
rect 9956 11160 10008 11212
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 4896 11092 4948 11144
rect 5816 11092 5868 11144
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 6368 11024 6420 11076
rect 6736 11092 6788 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7288 11092 7340 11144
rect 4528 10956 4580 11008
rect 5908 10956 5960 11008
rect 6000 10956 6052 11008
rect 8300 11024 8352 11076
rect 8484 11024 8536 11076
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10784 11092 10836 11144
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11336 11092 11388 11144
rect 12348 11228 12400 11280
rect 9312 10956 9364 11008
rect 11428 11024 11480 11076
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 13544 11228 13596 11280
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 9772 10999 9824 11008
rect 9772 10965 9781 10999
rect 9781 10965 9815 10999
rect 9815 10965 9824 10999
rect 9772 10956 9824 10965
rect 9864 10956 9916 11008
rect 10692 10956 10744 11008
rect 11060 10956 11112 11008
rect 11888 10956 11940 11008
rect 12348 10956 12400 11008
rect 12532 10956 12584 11008
rect 4918 10854 4970 10906
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 5238 10854 5290 10906
rect 10918 10854 10970 10906
rect 10982 10854 11034 10906
rect 11046 10854 11098 10906
rect 11110 10854 11162 10906
rect 11174 10854 11226 10906
rect 11238 10854 11290 10906
rect 3424 10752 3476 10804
rect 3884 10752 3936 10804
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3332 10616 3384 10668
rect 4528 10684 4580 10736
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 3608 10548 3660 10600
rect 4068 10616 4120 10668
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 6000 10752 6052 10804
rect 7380 10752 7432 10804
rect 8392 10752 8444 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 9128 10752 9180 10804
rect 4160 10616 4212 10625
rect 5264 10616 5316 10668
rect 6736 10684 6788 10736
rect 5540 10616 5592 10668
rect 5632 10548 5684 10600
rect 3792 10523 3844 10532
rect 3792 10489 3801 10523
rect 3801 10489 3835 10523
rect 3835 10489 3844 10523
rect 3792 10480 3844 10489
rect 4804 10480 4856 10532
rect 6368 10616 6420 10668
rect 6644 10616 6696 10668
rect 7288 10616 7340 10668
rect 7564 10616 7616 10668
rect 7840 10616 7892 10668
rect 7196 10548 7248 10600
rect 7656 10548 7708 10600
rect 8116 10591 8168 10600
rect 8116 10557 8125 10591
rect 8125 10557 8159 10591
rect 8159 10557 8168 10591
rect 8116 10548 8168 10557
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 9680 10752 9732 10804
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 9956 10752 10008 10804
rect 10140 10752 10192 10804
rect 10324 10752 10376 10804
rect 10692 10752 10744 10804
rect 11336 10752 11388 10804
rect 11520 10752 11572 10804
rect 11612 10752 11664 10804
rect 11980 10752 12032 10804
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 8576 10548 8628 10600
rect 9588 10616 9640 10668
rect 10416 10684 10468 10736
rect 11244 10684 11296 10736
rect 9956 10616 10008 10668
rect 10048 10616 10100 10668
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10784 10616 10836 10668
rect 4528 10412 4580 10464
rect 6092 10480 6144 10532
rect 6184 10523 6236 10532
rect 6184 10489 6193 10523
rect 6193 10489 6227 10523
rect 6227 10489 6236 10523
rect 6184 10480 6236 10489
rect 6368 10480 6420 10532
rect 5448 10412 5500 10464
rect 6460 10412 6512 10464
rect 6552 10412 6604 10464
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 7196 10412 7248 10464
rect 7748 10480 7800 10532
rect 10508 10548 10560 10600
rect 12072 10616 12124 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12532 10548 12584 10600
rect 10048 10523 10100 10532
rect 10048 10489 10057 10523
rect 10057 10489 10091 10523
rect 10091 10489 10100 10523
rect 10048 10480 10100 10489
rect 12900 10548 12952 10600
rect 9220 10412 9272 10464
rect 9680 10412 9732 10464
rect 9864 10412 9916 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 12440 10412 12492 10464
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 2872 10208 2924 10260
rect 6184 10208 6236 10260
rect 7288 10208 7340 10260
rect 3424 10115 3476 10124
rect 3424 10081 3433 10115
rect 3433 10081 3467 10115
rect 3467 10081 3476 10115
rect 3424 10072 3476 10081
rect 7380 10072 7432 10124
rect 8392 10140 8444 10192
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 6552 10004 6604 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 3884 9936 3936 9988
rect 4344 9936 4396 9988
rect 4620 9936 4672 9988
rect 6828 9936 6880 9988
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 7656 10004 7708 10056
rect 7840 10004 7892 10056
rect 8300 10004 8352 10056
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 12164 10251 12216 10260
rect 12164 10217 12173 10251
rect 12173 10217 12207 10251
rect 12207 10217 12216 10251
rect 12164 10208 12216 10217
rect 9036 10004 9088 10056
rect 9220 10004 9272 10056
rect 9956 10140 10008 10192
rect 11428 10140 11480 10192
rect 12808 10140 12860 10192
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 9956 10004 10008 10056
rect 10140 10004 10192 10056
rect 2872 9868 2924 9920
rect 3332 9868 3384 9920
rect 3608 9868 3660 9920
rect 4160 9868 4212 9920
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 7012 9868 7064 9920
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 7564 9868 7616 9920
rect 8392 9868 8444 9920
rect 8484 9868 8536 9920
rect 9220 9911 9272 9920
rect 9220 9877 9229 9911
rect 9229 9877 9263 9911
rect 9263 9877 9272 9911
rect 9220 9868 9272 9877
rect 10508 9936 10560 9988
rect 10784 9936 10836 9988
rect 10600 9868 10652 9920
rect 11796 9868 11848 9920
rect 4918 9766 4970 9818
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 5238 9766 5290 9818
rect 10918 9766 10970 9818
rect 10982 9766 11034 9818
rect 11046 9766 11098 9818
rect 11110 9766 11162 9818
rect 11174 9766 11226 9818
rect 11238 9766 11290 9818
rect 3240 9707 3292 9716
rect 3240 9673 3249 9707
rect 3249 9673 3283 9707
rect 3283 9673 3292 9707
rect 3240 9664 3292 9673
rect 3976 9664 4028 9716
rect 3240 9528 3292 9580
rect 4896 9596 4948 9648
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 2872 9392 2924 9444
rect 1768 9324 1820 9376
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 3516 9460 3568 9512
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 3884 9460 3936 9512
rect 4528 9528 4580 9580
rect 4712 9528 4764 9580
rect 5816 9664 5868 9716
rect 7288 9664 7340 9716
rect 4252 9460 4304 9512
rect 5632 9528 5684 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6092 9596 6144 9648
rect 7012 9596 7064 9648
rect 8392 9664 8444 9716
rect 8576 9664 8628 9716
rect 10324 9664 10376 9716
rect 4896 9460 4948 9512
rect 6736 9528 6788 9580
rect 6644 9460 6696 9512
rect 5632 9392 5684 9444
rect 7012 9460 7064 9512
rect 6828 9392 6880 9444
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 8668 9596 8720 9648
rect 9220 9596 9272 9648
rect 10876 9664 10928 9716
rect 8484 9528 8536 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 8116 9460 8168 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 9588 9528 9640 9580
rect 10048 9528 10100 9580
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10416 9528 10468 9580
rect 11336 9596 11388 9648
rect 12072 9664 12124 9716
rect 12440 9596 12492 9648
rect 8760 9460 8812 9469
rect 8576 9392 8628 9444
rect 7104 9324 7156 9376
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 8944 9324 8996 9376
rect 9680 9324 9732 9376
rect 10692 9324 10744 9376
rect 10968 9561 11020 9580
rect 10968 9528 10978 9561
rect 10978 9528 11012 9561
rect 11012 9528 11020 9561
rect 10968 9392 11020 9444
rect 11520 9460 11572 9512
rect 12716 9392 12768 9444
rect 11704 9324 11756 9376
rect 12348 9324 12400 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 3424 9120 3476 9172
rect 4068 9120 4120 9172
rect 4344 9120 4396 9172
rect 2964 8984 3016 9036
rect 3424 8984 3476 9036
rect 3608 9027 3660 9036
rect 3608 8993 3617 9027
rect 3617 8993 3651 9027
rect 3651 8993 3660 9027
rect 3608 8984 3660 8993
rect 4436 9052 4488 9104
rect 4804 9120 4856 9172
rect 4896 9052 4948 9104
rect 2780 8916 2832 8968
rect 3056 8916 3108 8968
rect 3976 8916 4028 8968
rect 4252 8984 4304 9036
rect 1768 8891 1820 8900
rect 1768 8857 1802 8891
rect 1802 8857 1820 8891
rect 1768 8848 1820 8857
rect 4344 8916 4396 8968
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4712 8984 4764 9036
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3516 8823 3568 8832
rect 3516 8789 3525 8823
rect 3525 8789 3559 8823
rect 3559 8789 3568 8823
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5540 9120 5592 9172
rect 6644 9120 6696 9172
rect 7104 9120 7156 9172
rect 7380 9120 7432 9172
rect 5632 9052 5684 9104
rect 5448 8916 5500 8968
rect 5816 8984 5868 9036
rect 6368 8984 6420 9036
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 7656 9052 7708 9104
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7012 8984 7064 9036
rect 8944 9120 8996 9172
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 10324 9120 10376 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11060 9120 11112 9172
rect 11520 9120 11572 9172
rect 8852 9052 8904 9104
rect 9680 9052 9732 9104
rect 10140 9052 10192 9104
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 4712 8848 4764 8900
rect 7104 8891 7156 8900
rect 7104 8857 7113 8891
rect 7113 8857 7147 8891
rect 7147 8857 7156 8891
rect 7564 8916 7616 8968
rect 7656 8916 7708 8968
rect 7840 8916 7892 8968
rect 10324 8984 10376 9036
rect 10692 8984 10744 9036
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9312 8916 9364 8968
rect 9588 8916 9640 8968
rect 10876 8916 10928 8968
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 7104 8848 7156 8857
rect 8392 8848 8444 8900
rect 9864 8848 9916 8900
rect 10048 8848 10100 8900
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11428 8916 11480 8968
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 11980 8891 12032 8900
rect 11980 8857 11989 8891
rect 11989 8857 12023 8891
rect 12023 8857 12032 8891
rect 11980 8848 12032 8857
rect 3516 8780 3568 8789
rect 4620 8780 4672 8832
rect 4988 8780 5040 8832
rect 5448 8780 5500 8832
rect 7012 8780 7064 8832
rect 8484 8780 8536 8832
rect 10140 8780 10192 8832
rect 10416 8780 10468 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 4918 8678 4970 8730
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 5238 8678 5290 8730
rect 10918 8678 10970 8730
rect 10982 8678 11034 8730
rect 11046 8678 11098 8730
rect 11110 8678 11162 8730
rect 11174 8678 11226 8730
rect 11238 8678 11290 8730
rect 2964 8576 3016 8628
rect 3792 8576 3844 8628
rect 4252 8619 4304 8628
rect 4252 8585 4261 8619
rect 4261 8585 4295 8619
rect 4295 8585 4304 8619
rect 4252 8576 4304 8585
rect 4344 8576 4396 8628
rect 4528 8576 4580 8628
rect 5448 8576 5500 8628
rect 5816 8576 5868 8628
rect 6920 8576 6972 8628
rect 10508 8576 10560 8628
rect 4068 8508 4120 8560
rect 3976 8440 4028 8492
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 7288 8508 7340 8560
rect 14188 8508 14240 8560
rect 10784 8440 10836 8492
rect 12440 8440 12492 8492
rect 13544 8440 13596 8492
rect 3424 8304 3476 8356
rect 3700 8304 3752 8356
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 5908 8372 5960 8424
rect 6368 8372 6420 8424
rect 7656 8372 7708 8424
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 4712 8236 4764 8288
rect 4896 8236 4948 8288
rect 8392 8304 8444 8356
rect 9128 8304 9180 8356
rect 7012 8279 7064 8288
rect 7012 8245 7021 8279
rect 7021 8245 7055 8279
rect 7055 8245 7064 8279
rect 7012 8236 7064 8245
rect 9496 8236 9548 8288
rect 12164 8236 12216 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 5632 8032 5684 8084
rect 6828 8032 6880 8084
rect 7840 8032 7892 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 10048 8032 10100 8084
rect 10600 8032 10652 8084
rect 11980 8032 12032 8084
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 4620 7828 4672 7880
rect 9588 7896 9640 7948
rect 11520 7896 11572 7948
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 5724 7828 5776 7880
rect 7840 7828 7892 7880
rect 8944 7828 8996 7880
rect 9036 7760 9088 7812
rect 9312 7803 9364 7812
rect 9312 7769 9321 7803
rect 9321 7769 9355 7803
rect 9355 7769 9364 7803
rect 9312 7760 9364 7769
rect 9864 7828 9916 7880
rect 10324 7828 10376 7880
rect 10784 7828 10836 7880
rect 2596 7735 2648 7744
rect 2596 7701 2605 7735
rect 2605 7701 2639 7735
rect 2639 7701 2648 7735
rect 2596 7692 2648 7701
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10600 7760 10652 7812
rect 11796 7828 11848 7880
rect 12072 7828 12124 7880
rect 12900 7896 12952 7948
rect 12440 7871 12492 7880
rect 12440 7837 12449 7871
rect 12449 7837 12483 7871
rect 12483 7837 12492 7871
rect 12440 7828 12492 7837
rect 12808 7760 12860 7812
rect 11336 7692 11388 7744
rect 12532 7692 12584 7744
rect 4918 7590 4970 7642
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 5238 7590 5290 7642
rect 10918 7590 10970 7642
rect 10982 7590 11034 7642
rect 11046 7590 11098 7642
rect 11110 7590 11162 7642
rect 11174 7590 11226 7642
rect 11238 7590 11290 7642
rect 2596 7488 2648 7540
rect 3792 7488 3844 7540
rect 9036 7531 9088 7540
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 10232 7488 10284 7540
rect 11060 7488 11112 7540
rect 11428 7488 11480 7540
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 8300 7352 8352 7404
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 8760 7352 8812 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 9864 7420 9916 7472
rect 9680 7352 9732 7404
rect 3884 7216 3936 7268
rect 7748 7216 7800 7268
rect 8760 7216 8812 7268
rect 10600 7352 10652 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 12808 7352 12860 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 2412 7148 2464 7200
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4712 7148 4764 7200
rect 6092 7148 6144 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7288 7148 7340 7200
rect 9772 7148 9824 7200
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 10876 7148 10928 7200
rect 11980 7148 12032 7200
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 4252 6944 4304 6996
rect 5724 6944 5776 6996
rect 7840 6944 7892 6996
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 9404 6944 9456 6996
rect 10232 6944 10284 6996
rect 10324 6944 10376 6996
rect 10876 6944 10928 6996
rect 8944 6876 8996 6928
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4344 6783 4396 6792
rect 4344 6749 4378 6783
rect 4378 6749 4396 6783
rect 4344 6740 4396 6749
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 7196 6740 7248 6792
rect 7932 6740 7984 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 8392 6672 8444 6724
rect 8668 6672 8720 6724
rect 9220 6672 9272 6724
rect 10600 6876 10652 6928
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10692 6740 10744 6792
rect 11796 6944 11848 6996
rect 11152 6876 11204 6928
rect 11428 6876 11480 6928
rect 11428 6783 11480 6786
rect 11428 6749 11444 6783
rect 11444 6749 11478 6783
rect 11478 6749 11480 6783
rect 11428 6734 11480 6749
rect 11980 6740 12032 6792
rect 12072 6740 12124 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 4918 6502 4970 6554
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 5238 6502 5290 6554
rect 10918 6502 10970 6554
rect 10982 6502 11034 6554
rect 11046 6502 11098 6554
rect 11110 6502 11162 6554
rect 11174 6502 11226 6554
rect 11238 6502 11290 6554
rect 4436 6400 4488 6452
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2872 6332 2924 6384
rect 3516 6332 3568 6384
rect 6920 6332 6972 6384
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 3608 6264 3660 6316
rect 7196 6400 7248 6452
rect 7288 6400 7340 6452
rect 7104 6332 7156 6384
rect 7748 6332 7800 6384
rect 8576 6400 8628 6452
rect 8760 6400 8812 6452
rect 8852 6400 8904 6452
rect 2596 6196 2648 6248
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7564 6307 7616 6316
rect 7564 6273 7572 6307
rect 7572 6273 7606 6307
rect 7606 6273 7616 6307
rect 7564 6264 7616 6273
rect 7012 6196 7064 6248
rect 8484 6264 8536 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 9220 6332 9272 6384
rect 9680 6332 9732 6384
rect 9772 6332 9824 6384
rect 9956 6332 10008 6384
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 10324 6264 10376 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 4068 6128 4120 6180
rect 1768 6060 1820 6112
rect 2780 6060 2832 6112
rect 6644 6171 6696 6180
rect 6644 6137 6653 6171
rect 6653 6137 6687 6171
rect 6687 6137 6696 6171
rect 6644 6128 6696 6137
rect 7748 6128 7800 6180
rect 8392 6128 8444 6180
rect 9496 6196 9548 6248
rect 10140 6196 10192 6248
rect 11336 6400 11388 6452
rect 11060 6264 11112 6316
rect 11520 6264 11572 6316
rect 11888 6264 11940 6316
rect 12900 6264 12952 6316
rect 10048 6128 10100 6180
rect 6184 6060 6236 6112
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 7564 6060 7616 6112
rect 8852 6060 8904 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 9220 6103 9272 6112
rect 9220 6069 9229 6103
rect 9229 6069 9263 6103
rect 9263 6069 9272 6103
rect 9220 6060 9272 6069
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 12808 6196 12860 6248
rect 11428 6128 11480 6180
rect 11336 6060 11388 6112
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 2504 5856 2556 5908
rect 4160 5788 4212 5840
rect 1768 5584 1820 5636
rect 4068 5652 4120 5704
rect 4804 5652 4856 5704
rect 6184 5856 6236 5908
rect 7012 5856 7064 5908
rect 2780 5516 2832 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 4344 5584 4396 5636
rect 7196 5652 7248 5704
rect 7748 5652 7800 5704
rect 6644 5584 6696 5636
rect 9496 5856 9548 5908
rect 9864 5856 9916 5908
rect 10324 5856 10376 5908
rect 8576 5788 8628 5840
rect 8760 5788 8812 5840
rect 9404 5788 9456 5840
rect 10600 5788 10652 5840
rect 11704 5788 11756 5840
rect 9036 5652 9088 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10324 5652 10376 5704
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 7380 5516 7432 5568
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 9864 5516 9916 5568
rect 11244 5516 11296 5568
rect 11520 5516 11572 5568
rect 4918 5414 4970 5466
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 5238 5414 5290 5466
rect 10918 5414 10970 5466
rect 10982 5414 11034 5466
rect 11046 5414 11098 5466
rect 11110 5414 11162 5466
rect 11174 5414 11226 5466
rect 11238 5414 11290 5466
rect 2872 5312 2924 5364
rect 2780 5176 2832 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3792 5312 3844 5364
rect 4068 5312 4120 5364
rect 7104 5312 7156 5364
rect 9128 5312 9180 5364
rect 10232 5312 10284 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3792 5176 3844 5228
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4804 5176 4856 5228
rect 5448 5176 5500 5228
rect 6920 5176 6972 5228
rect 9036 5176 9088 5228
rect 9404 5176 9456 5228
rect 4068 5108 4120 5160
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 10324 5176 10376 5228
rect 10416 5176 10468 5228
rect 11336 5176 11388 5228
rect 11428 5176 11480 5228
rect 1584 4972 1636 5024
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4160 4972 4212 5024
rect 5540 4972 5592 5024
rect 10232 4972 10284 5024
rect 11336 4972 11388 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 4068 4768 4120 4820
rect 8576 4768 8628 4820
rect 8944 4768 8996 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 3792 4564 3844 4616
rect 4528 4564 4580 4616
rect 4712 4564 4764 4616
rect 5540 4632 5592 4684
rect 4620 4496 4672 4548
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 8852 4564 8904 4616
rect 10416 4768 10468 4820
rect 10232 4700 10284 4752
rect 6368 4496 6420 4548
rect 9680 4496 9732 4548
rect 9956 4564 10008 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10324 4632 10376 4684
rect 11520 4632 11572 4684
rect 11796 4564 11848 4616
rect 4712 4471 4764 4480
rect 4712 4437 4721 4471
rect 4721 4437 4755 4471
rect 4755 4437 4764 4471
rect 4712 4428 4764 4437
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 8392 4428 8444 4480
rect 9220 4428 9272 4480
rect 9588 4428 9640 4480
rect 10692 4428 10744 4480
rect 13452 4496 13504 4548
rect 4918 4326 4970 4378
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 5238 4326 5290 4378
rect 10918 4326 10970 4378
rect 10982 4326 11034 4378
rect 11046 4326 11098 4378
rect 11110 4326 11162 4378
rect 11174 4326 11226 4378
rect 11238 4326 11290 4378
rect 2872 4224 2924 4276
rect 3700 4224 3752 4276
rect 5540 4224 5592 4276
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 7104 4224 7156 4276
rect 2780 4088 2832 4140
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 3976 4156 4028 4208
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 3516 4063 3568 4072
rect 3516 4029 3525 4063
rect 3525 4029 3559 4063
rect 3559 4029 3568 4063
rect 3516 4020 3568 4029
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 6644 4088 6696 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 8576 4224 8628 4276
rect 6828 4088 6880 4097
rect 7288 4088 7340 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 9680 4224 9732 4276
rect 13452 4224 13504 4276
rect 9956 4156 10008 4208
rect 11520 4156 11572 4208
rect 8392 4088 8444 4140
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 2596 3884 2648 3936
rect 4252 3884 4304 3936
rect 6184 3884 6236 3936
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 8944 4088 8996 4140
rect 9220 4088 9272 4140
rect 9772 4088 9824 4140
rect 13544 4088 13596 4140
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 8944 3884 8996 3936
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12072 3884 12124 3936
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 4436 3680 4488 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 12164 3680 12216 3732
rect 7288 3612 7340 3664
rect 3516 3544 3568 3596
rect 4068 3544 4120 3596
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4252 3476 4304 3528
rect 6184 3519 6236 3528
rect 6184 3485 6218 3519
rect 6218 3485 6236 3519
rect 6184 3476 6236 3485
rect 9956 3476 10008 3528
rect 10692 3519 10744 3528
rect 10692 3485 10726 3519
rect 10726 3485 10744 3519
rect 10692 3476 10744 3485
rect 2596 3408 2648 3460
rect 4804 3408 4856 3460
rect 7748 3408 7800 3460
rect 8668 3408 8720 3460
rect 8852 3408 8904 3460
rect 9036 3408 9088 3460
rect 3608 3383 3660 3392
rect 3608 3349 3617 3383
rect 3617 3349 3651 3383
rect 3651 3349 3660 3383
rect 3608 3340 3660 3349
rect 7564 3340 7616 3392
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 4918 3238 4970 3290
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 5238 3238 5290 3290
rect 10918 3238 10970 3290
rect 10982 3238 11034 3290
rect 11046 3238 11098 3290
rect 11110 3238 11162 3290
rect 11174 3238 11226 3290
rect 11238 3238 11290 3290
rect 3240 3136 3292 3188
rect 3608 3136 3660 3188
rect 5632 3136 5684 3188
rect 7564 3136 7616 3188
rect 8668 3179 8720 3188
rect 8668 3145 8677 3179
rect 8677 3145 8711 3179
rect 8711 3145 8720 3179
rect 8668 3136 8720 3145
rect 8760 3136 8812 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 10324 3136 10376 3188
rect 4160 3068 4212 3120
rect 4712 3068 4764 3120
rect 6828 3068 6880 3120
rect 8576 3068 8628 3120
rect 3884 3000 3936 3052
rect 4068 3000 4120 3052
rect 6644 3000 6696 3052
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 6000 2839 6052 2848
rect 6000 2805 6009 2839
rect 6009 2805 6043 2839
rect 6043 2805 6052 2839
rect 6000 2796 6052 2805
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 4620 2592 4672 2644
rect 6644 2592 6696 2644
rect 13544 2635 13596 2644
rect 13544 2601 13553 2635
rect 13553 2601 13587 2635
rect 13587 2601 13596 2635
rect 13544 2592 13596 2601
rect 4160 2524 4212 2576
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2964 2388 3016 2440
rect 3424 2388 3476 2440
rect 4252 2388 4304 2440
rect 6000 2456 6052 2508
rect 6828 2388 6880 2440
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7564 2388 7616 2440
rect 9864 2388 9916 2440
rect 10416 2388 10468 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12164 2388 12216 2440
rect 14188 2388 14240 2440
rect 1032 2252 1084 2304
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 3424 2252 3476 2304
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 5908 2295 5960 2304
rect 5908 2261 5917 2295
rect 5917 2261 5951 2295
rect 5951 2261 5960 2295
rect 5908 2252 5960 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 8208 2252 8260 2304
rect 9496 2295 9548 2304
rect 9496 2261 9505 2295
rect 9505 2261 9539 2295
rect 9539 2261 9548 2295
rect 9496 2252 9548 2261
rect 10692 2295 10744 2304
rect 10692 2261 10701 2295
rect 10701 2261 10735 2295
rect 10735 2261 10744 2295
rect 10692 2252 10744 2261
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 4918 2150 4970 2202
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 5238 2150 5290 2202
rect 10918 2150 10970 2202
rect 10982 2150 11034 2202
rect 11046 2150 11098 2202
rect 11110 2150 11162 2202
rect 11174 2150 11226 2202
rect 11238 2150 11290 2202
<< metal2 >>
rect 1030 16589 1086 17389
rect 2042 16589 2098 17389
rect 2148 16646 2360 16674
rect 1044 14618 1072 16589
rect 2056 16538 2084 16589
rect 2148 16538 2176 16646
rect 2056 16510 2176 16538
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2332 14618 2360 16646
rect 3054 16589 3110 17389
rect 4066 16589 4122 17389
rect 5078 16589 5134 17389
rect 6090 16589 6146 17389
rect 7102 16589 7158 17389
rect 7852 16646 8064 16674
rect 3068 14618 3096 16589
rect 4080 14618 4108 16589
rect 5092 14618 5120 16589
rect 6104 14618 6132 16589
rect 7116 14618 7144 16589
rect 7852 14618 7880 16646
rect 8036 16538 8064 16646
rect 8114 16589 8170 17389
rect 9126 16589 9182 17389
rect 10138 16589 10194 17389
rect 11150 16589 11206 17389
rect 12162 16589 12218 17389
rect 13174 16589 13230 17389
rect 14186 16589 14242 17389
rect 8128 16538 8156 16589
rect 8036 16510 8156 16538
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 9140 14618 9168 16589
rect 1032 14612 1084 14618
rect 1032 14554 1084 14560
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2148 12918 2176 13262
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2332 12986 2360 13194
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2228 12844 2280 12850
rect 2280 12804 2360 12832
rect 2228 12786 2280 12792
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 2332 12442 2360 12804
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 2516 11354 2544 14350
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2884 11218 2912 13262
rect 2976 12850 3004 13670
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12434 3372 12582
rect 3252 12406 3372 12434
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2976 11898 3004 12106
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 2884 10266 2912 11154
rect 2976 10606 3004 11494
rect 3068 10606 3096 11630
rect 3252 11121 3280 12406
rect 3436 12374 3464 13466
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3436 11257 3464 12310
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 3332 11144 3384 11150
rect 3238 11112 3294 11121
rect 3332 11086 3384 11092
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3238 11047 3294 11056
rect 3344 10674 3372 11086
rect 3436 10810 3464 11086
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3148 10668 3200 10674
rect 3332 10668 3384 10674
rect 3200 10628 3280 10656
rect 3148 10610 3200 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2872 10260 2924 10266
rect 2792 10220 2872 10248
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 8906 1808 9318
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 2318 9072 2374 9081
rect 2318 9007 2374 9016
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2332 6322 2360 9007
rect 2792 8974 2820 10220
rect 2872 10202 2924 10208
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9450 2912 9862
rect 2976 9518 3004 10542
rect 3068 9518 3096 10542
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3252 10044 3280 10628
rect 3332 10610 3384 10616
rect 3424 10124 3476 10130
rect 3528 10112 3556 14350
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3712 12442 3740 13806
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13258 4200 13670
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 3988 12838 4200 12866
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3804 12306 3832 12582
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3988 12238 4016 12838
rect 4172 12782 4200 12838
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4080 12238 4108 12718
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4252 12232 4304 12238
rect 4068 12174 4120 12180
rect 4250 12200 4252 12209
rect 4304 12200 4306 12209
rect 3620 11898 3648 12174
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3608 11688 3660 11694
rect 3712 11676 3740 12038
rect 3896 11694 3924 12174
rect 4080 11762 4108 12174
rect 4250 12135 4306 12144
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3660 11648 3740 11676
rect 3884 11688 3936 11694
rect 3608 11630 3660 11636
rect 3884 11630 3936 11636
rect 3620 10606 3648 11630
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3476 10084 3556 10112
rect 3424 10066 3476 10072
rect 3332 10056 3384 10062
rect 3252 10016 3332 10044
rect 3160 9568 3188 9998
rect 3252 9722 3280 10016
rect 3332 9998 3384 10004
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3240 9580 3292 9586
rect 3160 9540 3240 9568
rect 3240 9522 3292 9528
rect 3344 9518 3372 9862
rect 3528 9738 3556 10084
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3436 9710 3556 9738
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2976 9042 3004 9454
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3068 8974 3096 9454
rect 3436 9178 3464 9710
rect 3620 9625 3648 9862
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8634 3004 8774
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3436 8362 3464 8978
rect 3528 8838 3556 9454
rect 3620 9042 3648 9551
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3712 8362 3740 11154
rect 3896 10810 3924 11630
rect 4264 11354 4292 12135
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3988 10764 4200 10792
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3804 10169 3832 10474
rect 3790 10160 3846 10169
rect 3790 10095 3846 10104
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3896 9518 3924 9930
rect 3988 9722 4016 10764
rect 4172 10674 4200 10764
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4080 9908 4108 10610
rect 4160 9920 4212 9926
rect 4080 9880 4160 9908
rect 4160 9862 4212 9868
rect 4264 9738 4292 11086
rect 4356 9994 4384 14350
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4172 9710 4292 9738
rect 4172 9674 4200 9710
rect 4172 9646 4292 9674
rect 4264 9602 4292 9646
rect 4172 9574 4292 9602
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3804 8634 3832 9454
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 2792 7886 2820 8230
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7546 2636 7686
rect 3804 7546 3832 8230
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3896 7274 3924 9454
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8498 4016 8910
rect 4080 8566 4108 9114
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 2424 6914 2452 7142
rect 2424 6886 2636 6914
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5642 1808 6054
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 2516 5914 2544 6258
rect 2608 6254 2636 6886
rect 3528 6390 3556 7142
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 2792 5574 2820 6054
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5234 2820 5510
rect 2884 5370 2912 6326
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 3238 5536 3294 5545
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 2446 1624 4966
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 2792 4146 2820 5170
rect 2884 4282 2912 5306
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 2608 3466 2636 3878
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 2976 2446 3004 5510
rect 3238 5471 3294 5480
rect 3252 5234 3280 5471
rect 3620 5234 3648 6258
rect 4080 6186 4108 6802
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4172 5846 4200 9574
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 9042 4292 9454
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8634 4292 8978
rect 4356 8974 4384 9114
rect 4448 9110 4476 14350
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 4916 14172 5292 14181
rect 4972 14170 4996 14172
rect 5052 14170 5076 14172
rect 5132 14170 5156 14172
rect 5212 14170 5236 14172
rect 4972 14118 4982 14170
rect 5226 14118 5236 14170
rect 4972 14116 4996 14118
rect 5052 14116 5076 14118
rect 5132 14116 5156 14118
rect 5212 14116 5236 14118
rect 4916 14107 5292 14116
rect 5460 13938 5488 14282
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 4540 12442 4568 13738
rect 5276 13530 5304 13738
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4988 13456 5040 13462
rect 4816 13416 4988 13444
rect 4816 12782 4844 13416
rect 4988 13398 5040 13404
rect 4916 13084 5292 13093
rect 4972 13082 4996 13084
rect 5052 13082 5076 13084
rect 5132 13082 5156 13084
rect 5212 13082 5236 13084
rect 4972 13030 4982 13082
rect 5226 13030 5236 13082
rect 4972 13028 4996 13030
rect 5052 13028 5076 13030
rect 5132 13028 5156 13030
rect 5212 13028 5236 13030
rect 4916 13019 5292 13028
rect 5368 12986 5396 13874
rect 5460 13530 5488 13874
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4908 12782 4936 12854
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11898 4568 12174
rect 4632 12102 4660 12650
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4528 11892 4580 11898
rect 4816 11880 4844 12718
rect 4908 12374 4936 12718
rect 5184 12442 5212 12718
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4908 12102 4936 12174
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4916 11996 5292 12005
rect 4972 11994 4996 11996
rect 5052 11994 5076 11996
rect 5132 11994 5156 11996
rect 5212 11994 5236 11996
rect 4972 11942 4982 11994
rect 5226 11942 5236 11994
rect 4972 11940 4996 11942
rect 5052 11940 5076 11942
rect 5132 11940 5156 11942
rect 5212 11940 5236 11942
rect 4916 11931 5292 11940
rect 4816 11852 5212 11880
rect 4528 11834 4580 11840
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10742 4568 10950
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4528 10464 4580 10470
rect 4632 10452 4660 11698
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4724 11082 4752 11494
rect 4908 11150 4936 11698
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4816 10656 4844 11086
rect 5184 10996 5212 11852
rect 5368 11286 5396 12310
rect 5460 12306 5488 13126
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 12170 5580 12242
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5184 10968 5396 10996
rect 4916 10908 5292 10917
rect 4972 10906 4996 10908
rect 5052 10906 5076 10908
rect 5132 10906 5156 10908
rect 5212 10906 5236 10908
rect 4972 10854 4982 10906
rect 5226 10854 5236 10906
rect 4972 10852 4996 10854
rect 5052 10852 5076 10854
rect 5132 10852 5156 10854
rect 5212 10852 5236 10854
rect 4916 10843 5292 10852
rect 5368 10792 5396 10968
rect 4580 10424 4660 10452
rect 4724 10628 4844 10656
rect 5184 10764 5396 10792
rect 4528 10406 4580 10412
rect 4540 9586 4568 10406
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9364 4568 9522
rect 4632 9489 4660 9930
rect 4724 9586 4752 10628
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4618 9480 4674 9489
rect 4674 9438 4752 9466
rect 4618 9415 4674 9424
rect 4540 9336 4660 9364
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8634 4384 8910
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 5370 3832 5510
rect 4080 5370 4108 5646
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3792 5364 3844 5370
rect 4068 5364 4120 5370
rect 3792 5306 3844 5312
rect 3896 5324 4068 5352
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4622 3832 5170
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4298 3832 4558
rect 3712 4282 3832 4298
rect 3700 4276 3832 4282
rect 3752 4270 3832 4276
rect 3700 4218 3752 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3068 4049 3096 4082
rect 3054 4040 3110 4049
rect 3054 3975 3110 3984
rect 3252 3194 3280 4082
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3528 3602 3556 4014
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3896 3534 3924 5324
rect 4068 5306 4120 5312
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4214 4016 4966
rect 4080 4826 4108 5102
rect 4172 5030 4200 5510
rect 4264 5234 4292 6938
rect 4356 6798 4384 7686
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4448 6458 4476 9046
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8634 4568 8910
rect 4632 8838 4660 9336
rect 4724 9042 4752 9438
rect 4816 9178 4844 10474
rect 5184 9908 5212 10764
rect 5552 10674 5580 12106
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5276 10033 5304 10610
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5262 10024 5318 10033
rect 5262 9959 5318 9968
rect 5184 9880 5396 9908
rect 4916 9820 5292 9829
rect 4972 9818 4996 9820
rect 5052 9818 5076 9820
rect 5132 9818 5156 9820
rect 5212 9818 5236 9820
rect 4972 9766 4982 9818
rect 5226 9766 5236 9818
rect 4972 9764 4996 9766
rect 5052 9764 5076 9766
rect 5132 9764 5156 9766
rect 5212 9764 5236 9766
rect 4916 9755 5292 9764
rect 5368 9704 5396 9880
rect 5092 9676 5396 9704
rect 4896 9648 4948 9654
rect 4894 9616 4896 9625
rect 4948 9616 4950 9625
rect 4894 9551 4950 9560
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 9110 4936 9454
rect 4896 9104 4948 9110
rect 5092 9081 5120 9676
rect 4896 9046 4948 9052
rect 5078 9072 5134 9081
rect 4712 9036 4764 9042
rect 4764 8996 4844 9024
rect 5078 9007 5134 9016
rect 4712 8978 4764 8984
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4540 8498 4568 8570
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4724 8378 4752 8842
rect 4816 8498 4844 8996
rect 5460 8974 5488 10406
rect 5552 9178 5580 10610
rect 5632 10600 5684 10606
rect 5630 10568 5632 10577
rect 5684 10568 5686 10577
rect 5630 10503 5686 10512
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5644 9450 5672 9522
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 4896 8968 4948 8974
rect 5448 8968 5500 8974
rect 4948 8945 5028 8956
rect 4948 8936 5042 8945
rect 4948 8928 4986 8936
rect 4896 8910 4948 8916
rect 5448 8910 5500 8916
rect 4986 8871 5042 8880
rect 5000 8838 5028 8871
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4916 8732 5292 8741
rect 4972 8730 4996 8732
rect 5052 8730 5076 8732
rect 5132 8730 5156 8732
rect 5212 8730 5236 8732
rect 4972 8678 4982 8730
rect 5226 8678 5236 8730
rect 4972 8676 4996 8678
rect 5052 8676 5076 8678
rect 5132 8676 5156 8678
rect 5212 8676 5236 8678
rect 4916 8667 5292 8676
rect 5460 8634 5488 8774
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4896 8424 4948 8430
rect 4724 8372 4896 8378
rect 4724 8366 4948 8372
rect 4724 8350 4936 8366
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4712 8288 4764 8294
rect 4896 8288 4948 8294
rect 4764 8248 4896 8276
rect 4712 8230 4764 8236
rect 4896 8230 4948 8236
rect 4632 7886 4660 8230
rect 5644 8090 5672 9046
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 7886 5764 14350
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13258 6408 13670
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12442 6592 12786
rect 6748 12442 6776 13874
rect 6840 12646 6868 13874
rect 6932 13190 6960 14350
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7024 12850 7052 13874
rect 7116 12986 7144 13874
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 12986 7236 13670
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7300 12850 7328 13874
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 8404 13530 8432 14350
rect 9416 13734 9444 14350
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9692 13530 9720 13874
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 7668 12986 7696 13194
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 8312 12850 8340 13194
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7012 12844 7064 12850
rect 7288 12844 7340 12850
rect 7064 12804 7144 12832
rect 7012 12786 7064 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6932 12374 6960 12786
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 7024 12238 7052 12650
rect 7116 12434 7144 12804
rect 7288 12786 7340 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7116 12406 7512 12434
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 5828 11830 5856 12174
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 7024 11762 7052 12038
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 9722 5856 11086
rect 6380 11082 6408 11698
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9042 5856 9522
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 4916 7644 5292 7653
rect 4972 7642 4996 7644
rect 5052 7642 5076 7644
rect 5132 7642 5156 7644
rect 5212 7642 5236 7644
rect 4972 7590 4982 7642
rect 5226 7590 5236 7642
rect 4972 7588 4996 7590
rect 5052 7588 5076 7590
rect 5132 7588 5156 7590
rect 5212 7588 5236 7590
rect 4916 7579 5292 7588
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4356 5234 4384 5578
rect 4448 5386 4476 6394
rect 4448 5358 4568 5386
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3620 3194 3648 3334
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3620 2774 3648 3130
rect 3896 3058 3924 3470
rect 4080 3058 4108 3538
rect 4264 3534 4292 3878
rect 4448 3738 4476 5170
rect 4540 4622 4568 5358
rect 4724 4622 4752 7142
rect 5736 7002 5764 7822
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 4916 6556 5292 6565
rect 4972 6554 4996 6556
rect 5052 6554 5076 6556
rect 5132 6554 5156 6556
rect 5212 6554 5236 6556
rect 4972 6502 4982 6554
rect 5226 6502 5236 6554
rect 4972 6500 4996 6502
rect 5052 6500 5076 6502
rect 5132 6500 5156 6502
rect 5212 6500 5236 6502
rect 4916 6491 5292 6500
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5234 4844 5646
rect 4916 5468 5292 5477
rect 4972 5466 4996 5468
rect 5052 5466 5076 5468
rect 5132 5466 5156 5468
rect 5212 5466 5236 5468
rect 4972 5414 4982 5466
rect 5226 5414 5236 5466
rect 4972 5412 4996 5414
rect 5052 5412 5076 5414
rect 5132 5412 5156 5414
rect 5212 5412 5236 5414
rect 4916 5403 5292 5412
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4622 5488 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4690 5580 4966
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4172 3126 4200 3470
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3436 2746 3648 2774
rect 3436 2446 3464 2746
rect 4172 2582 4200 3062
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4264 2446 4292 3470
rect 4632 2650 4660 4490
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4724 3126 4752 4422
rect 4816 3466 4844 4422
rect 4916 4380 5292 4389
rect 4972 4378 4996 4380
rect 5052 4378 5076 4380
rect 5132 4378 5156 4380
rect 5212 4378 5236 4380
rect 4972 4326 4982 4378
rect 5226 4326 5236 4378
rect 4972 4324 4996 4326
rect 5052 4324 5076 4326
rect 5132 4324 5156 4326
rect 5212 4324 5236 4326
rect 4916 4315 5292 4324
rect 5460 4146 5488 4558
rect 5552 4282 5580 4626
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5828 4146 5856 8570
rect 5920 8430 5948 10950
rect 6012 10810 6040 10950
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 8974 6040 10746
rect 6380 10674 6408 11018
rect 6748 10742 6776 11086
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6368 10668 6420 10674
rect 6644 10668 6696 10674
rect 6368 10610 6420 10616
rect 6564 10628 6644 10656
rect 6380 10538 6408 10610
rect 6564 10588 6592 10628
rect 6644 10610 6696 10616
rect 6472 10560 6592 10588
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6104 9654 6132 10474
rect 6196 10266 6224 10474
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6380 9042 6408 10474
rect 6472 10470 6500 10560
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10062 6592 10406
rect 7024 10282 7052 11698
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 10470 7144 11630
rect 7300 11150 7328 12106
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11558 7420 11698
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 11354 7420 11494
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7208 10606 7236 11086
rect 7300 10674 7328 11086
rect 7392 10810 7420 11290
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7378 10704 7434 10713
rect 7288 10668 7340 10674
rect 7378 10639 7434 10648
rect 7288 10610 7340 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7024 10254 7144 10282
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9518 6684 9998
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6840 9874 6868 9930
rect 7012 9920 7064 9926
rect 6748 9586 6776 9862
rect 6840 9846 6960 9874
rect 7012 9862 7064 9868
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 9178 6684 9454
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6748 9081 6776 9522
rect 6826 9480 6882 9489
rect 6826 9415 6828 9424
rect 6880 9415 6882 9424
rect 6828 9386 6880 9392
rect 6734 9072 6790 9081
rect 6368 9036 6420 9042
rect 6734 9007 6790 9016
rect 6368 8978 6420 8984
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6380 8430 6408 8978
rect 6840 8974 6868 9386
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 5920 6798 5948 8366
rect 6840 8090 6868 8910
rect 6932 8634 6960 9846
rect 7024 9654 7052 9862
rect 7116 9738 7144 10254
rect 7208 10062 7236 10406
rect 7300 10266 7328 10610
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7392 10130 7420 10639
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7194 9752 7250 9761
rect 7116 9710 7194 9738
rect 7300 9722 7328 9862
rect 7194 9687 7250 9696
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7012 9648 7064 9654
rect 7010 9616 7012 9625
rect 7064 9616 7066 9625
rect 7010 9551 7066 9560
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7024 9042 7052 9454
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 9178 7144 9318
rect 7392 9178 7420 9522
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8838 7052 8978
rect 7288 8968 7340 8974
rect 7102 8936 7158 8945
rect 7288 8910 7340 8916
rect 7102 8871 7104 8880
rect 7156 8871 7158 8880
rect 7104 8842 7156 8848
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6798 6132 7142
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6118 6224 6734
rect 6932 6390 6960 8570
rect 7300 8566 7328 8910
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7410 7052 8230
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7208 6798 7236 7142
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 6458 7236 6734
rect 7300 6458 7328 7142
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7012 6248 7064 6254
rect 7010 6216 7012 6225
rect 7064 6216 7066 6225
rect 6644 6180 6696 6186
rect 7010 6151 7066 6160
rect 6644 6122 6696 6128
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5914 6224 6054
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6656 5642 6684 6122
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5914 7052 6054
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4282 6408 4490
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6656 4146 6684 5578
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5234 6960 5510
rect 7116 5370 7144 6326
rect 7208 5710 7236 6394
rect 7288 6316 7340 6322
rect 7340 6276 7420 6304
rect 7288 6258 7340 6264
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7392 5574 7420 6276
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7116 4282 7144 5306
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4916 3292 5292 3301
rect 4972 3290 4996 3292
rect 5052 3290 5076 3292
rect 5132 3290 5156 3292
rect 5212 3290 5236 3292
rect 4972 3238 4982 3290
rect 5226 3238 5236 3290
rect 4972 3236 4996 3238
rect 5052 3236 5076 3238
rect 5132 3236 5156 3238
rect 5212 3236 5236 3238
rect 4916 3227 5292 3236
rect 5644 3194 5672 4082
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3534 6224 3878
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 6656 3058 6684 4082
rect 6840 3126 6868 4082
rect 7300 3670 7328 4082
rect 7484 3942 7512 12406
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 7668 12050 7696 12582
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 8404 12442 8432 12718
rect 8496 12646 8524 13466
rect 9784 13410 9812 13874
rect 10152 13705 10180 16589
rect 11164 14414 11192 16589
rect 12176 14414 12204 16589
rect 13188 14414 13216 16589
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 10916 14172 11292 14181
rect 10972 14170 10996 14172
rect 11052 14170 11076 14172
rect 11132 14170 11156 14172
rect 11212 14170 11236 14172
rect 10972 14118 10982 14170
rect 11226 14118 11236 14170
rect 10972 14116 10996 14118
rect 11052 14116 11076 14118
rect 11132 14116 11156 14118
rect 11212 14116 11236 14118
rect 10916 14107 11292 14116
rect 11532 13841 11560 14214
rect 12268 13841 12296 14214
rect 11518 13832 11574 13841
rect 10692 13796 10744 13802
rect 11518 13767 11574 13776
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 10692 13738 10744 13744
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9692 13382 9812 13410
rect 9692 13326 9720 13382
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12918 9260 13126
rect 9692 12986 9720 13262
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9968 12918 9996 13466
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9312 12912 9364 12918
rect 9864 12912 9916 12918
rect 9312 12854 9364 12860
rect 9862 12880 9864 12889
rect 9956 12912 10008 12918
rect 9916 12880 9918 12889
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8496 12238 8524 12582
rect 9140 12345 9168 12650
rect 9126 12336 9182 12345
rect 9126 12271 9182 12280
rect 9140 12238 9168 12271
rect 9232 12238 9260 12854
rect 9324 12782 9352 12854
rect 9956 12854 10008 12860
rect 9862 12815 9918 12824
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9876 12594 9904 12815
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 8116 12096 8168 12102
rect 7668 12022 7972 12050
rect 8116 12038 8168 12044
rect 7668 11898 7696 12022
rect 7944 11898 7972 12022
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8128 11694 8156 12038
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7838 10704 7894 10713
rect 7564 10668 7616 10674
rect 7838 10639 7840 10648
rect 7564 10610 7616 10616
rect 7892 10639 7894 10648
rect 7840 10610 7892 10616
rect 7576 9926 7604 10610
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10062 7696 10542
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7760 9674 7788 10474
rect 7944 10452 7972 11222
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8312 10674 8340 11018
rect 8496 10810 8524 11018
rect 9140 10810 9168 12174
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8116 10600 8168 10606
rect 8114 10568 8116 10577
rect 8168 10568 8170 10577
rect 8114 10503 8170 10512
rect 7852 10424 7972 10452
rect 7852 10146 7880 10424
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 8404 10198 8432 10746
rect 8576 10600 8628 10606
rect 8496 10560 8576 10588
rect 8392 10192 8444 10198
rect 8298 10160 8354 10169
rect 7852 10130 8156 10146
rect 7852 10124 8168 10130
rect 7852 10118 8116 10124
rect 8392 10134 8444 10140
rect 8298 10095 8354 10104
rect 8116 10066 8168 10072
rect 8312 10062 8340 10095
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7668 9646 7788 9674
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 8974 7604 9522
rect 7668 9110 7696 9646
rect 7656 9104 7708 9110
rect 7852 9058 7880 9998
rect 8496 9926 8524 10560
rect 8576 10542 8628 10548
rect 9232 10470 9260 12174
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8392 9920 8444 9926
rect 8390 9888 8392 9897
rect 8484 9920 8536 9926
rect 8444 9888 8446 9897
rect 8484 9862 8536 9868
rect 8390 9823 8446 9832
rect 8206 9752 8262 9761
rect 8206 9687 8262 9696
rect 8392 9716 8444 9722
rect 8116 9512 8168 9518
rect 8114 9480 8116 9489
rect 8168 9480 8170 9489
rect 8114 9415 8170 9424
rect 8116 9376 8168 9382
rect 8220 9364 8248 9687
rect 8392 9658 8444 9664
rect 8168 9336 8248 9364
rect 8116 9318 8168 9324
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 7656 9046 7708 9052
rect 7760 9030 7880 9058
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 8430 7696 8910
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7760 7274 7788 9030
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8090 7880 8910
rect 8404 8906 8432 9658
rect 8496 9586 8524 9862
rect 8588 9722 8616 10066
rect 9232 10062 9260 10406
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8668 9648 8720 9654
rect 8666 9616 8668 9625
rect 8720 9616 8722 9625
rect 8484 9580 8536 9586
rect 8666 9551 8722 9560
rect 8852 9580 8904 9586
rect 8484 9522 8536 9528
rect 8852 9522 8904 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8496 8838 8524 9522
rect 8760 9512 8812 9518
rect 8758 9480 8760 9489
rect 8812 9480 8814 9489
rect 8576 9444 8628 9450
rect 8758 9415 8814 9424
rect 8576 9386 8628 9392
rect 8588 9081 8616 9386
rect 8864 9110 8892 9522
rect 8956 9382 8984 9522
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9048 9178 9076 9998
rect 9220 9920 9272 9926
rect 9324 9897 9352 10950
rect 9416 10266 9444 11154
rect 9692 10810 9720 12582
rect 9876 12566 9996 12594
rect 9968 12356 9996 12566
rect 9876 12328 9996 12356
rect 9876 12238 9904 12328
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9784 11898 9812 12174
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11830 9904 12038
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10152 11880 10180 12242
rect 10244 12238 10272 13194
rect 10336 12442 10364 13262
rect 10704 13190 10732 13738
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12850 10732 13126
rect 10916 13084 11292 13093
rect 10972 13082 10996 13084
rect 11052 13082 11076 13084
rect 11132 13082 11156 13084
rect 11212 13082 11236 13084
rect 10972 13030 10982 13082
rect 11226 13030 11236 13082
rect 10972 13028 10996 13030
rect 11052 13028 11076 13030
rect 11132 13028 11156 13030
rect 11212 13028 11236 13030
rect 10916 13019 11292 13028
rect 11244 12980 11296 12986
rect 11164 12940 11244 12968
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10428 12152 10456 12378
rect 10336 12124 10456 12152
rect 10336 11914 10364 12124
rect 10520 12102 10548 12718
rect 10612 12238 10640 12786
rect 10704 12238 10732 12786
rect 10796 12646 10824 12786
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10508 12096 10560 12102
rect 10560 12044 10640 12050
rect 10508 12038 10640 12044
rect 10520 12022 10640 12038
rect 10336 11886 10456 11914
rect 10152 11852 10272 11880
rect 10048 11834 10100 11840
rect 9864 11824 9916 11830
rect 9770 11792 9826 11801
rect 9864 11766 9916 11772
rect 9770 11727 9772 11736
rect 9824 11727 9826 11736
rect 10048 11756 10100 11762
rect 9772 11698 9824 11704
rect 10048 11698 10100 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 11121 9996 11154
rect 9954 11112 10010 11121
rect 9954 11047 10010 11056
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 10690 9812 10950
rect 9876 10810 9904 10950
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9588 10668 9640 10674
rect 9784 10662 9904 10690
rect 9968 10674 9996 10746
rect 10060 10674 10088 11698
rect 10152 11150 10180 11698
rect 10244 11370 10272 11852
rect 10428 11694 10456 11886
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 11393 10548 11630
rect 10612 11626 10640 12022
rect 10704 11762 10732 12174
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10796 11694 10824 12310
rect 11164 12238 11192 12940
rect 11244 12922 11296 12928
rect 11348 12918 11376 13670
rect 12256 13252 12308 13258
rect 12176 13212 12256 13240
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12646 11376 12854
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11256 12434 11284 12582
rect 11256 12406 11376 12434
rect 11244 12368 11296 12374
rect 11242 12336 11244 12345
rect 11296 12336 11298 12345
rect 11242 12271 11298 12280
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10888 12102 10916 12174
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10916 11996 11292 12005
rect 10972 11994 10996 11996
rect 11052 11994 11076 11996
rect 11132 11994 11156 11996
rect 11212 11994 11236 11996
rect 10972 11942 10982 11994
rect 11226 11942 11236 11994
rect 10972 11940 10996 11942
rect 11052 11940 11076 11942
rect 11132 11940 11156 11942
rect 11212 11940 11236 11942
rect 10916 11931 11292 11940
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10506 11384 10562 11393
rect 10244 11342 10364 11370
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 11150 10272 11222
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10152 10810 10180 11086
rect 10336 10810 10364 11342
rect 10506 11319 10562 11328
rect 10414 11248 10470 11257
rect 10414 11183 10470 11192
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 9640 10628 9720 10656
rect 9588 10610 9640 10616
rect 9692 10588 9720 10628
rect 9692 10560 9812 10588
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9220 9862 9272 9868
rect 9310 9888 9366 9897
rect 9232 9654 9260 9862
rect 9310 9823 9366 9832
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8852 9104 8904 9110
rect 8574 9072 8630 9081
rect 8852 9046 8904 9052
rect 8574 9007 8630 9016
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 8404 7970 8432 8298
rect 8956 8090 8984 9114
rect 9324 8974 9352 9823
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 8974 9628 9522
rect 9692 9382 9720 10406
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9110 9720 9318
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9140 8362 9168 8910
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8312 7942 8432 7970
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 6390 7788 7210
rect 7852 7002 7880 7822
rect 8312 7410 8340 7942
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7932 6792 7984 6798
rect 8206 6760 8262 6769
rect 7984 6740 8206 6746
rect 7932 6734 8206 6740
rect 7944 6718 8206 6734
rect 7748 6384 7800 6390
rect 7944 6338 7972 6718
rect 8404 6730 8432 7686
rect 8956 7410 8984 7822
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9048 7546 9076 7754
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8760 7404 8812 7410
rect 8588 7364 8760 7392
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8496 7041 8524 7278
rect 8482 7032 8538 7041
rect 8482 6967 8538 6976
rect 8588 6798 8616 7364
rect 8760 7346 8812 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8772 6798 8800 7210
rect 9324 7002 9352 7754
rect 9402 7032 9458 7041
rect 9312 6996 9364 7002
rect 9402 6967 9404 6976
rect 9312 6938 9364 6944
rect 9456 6967 9458 6976
rect 9404 6938 9456 6944
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8206 6695 8262 6704
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8588 6458 8616 6734
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 7748 6326 7800 6332
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7852 6310 7972 6338
rect 8484 6316 8536 6322
rect 7576 6118 7604 6258
rect 7746 6216 7802 6225
rect 7746 6151 7748 6160
rect 7800 6151 7802 6160
rect 7748 6122 7800 6128
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7760 5710 7788 6122
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7852 4146 7880 6310
rect 8484 6258 8536 6264
rect 8392 6180 8444 6186
rect 8496 6168 8524 6258
rect 8444 6140 8524 6168
rect 8392 6122 8444 6128
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8588 5846 8616 6394
rect 8680 6322 8708 6666
rect 8772 6458 8800 6734
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8772 5846 8800 6394
rect 8864 6118 8892 6394
rect 8956 6322 8984 6870
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6390 9260 6666
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9324 6202 9352 6938
rect 9416 6322 9444 6938
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9508 6254 9536 8230
rect 9600 7954 9628 8910
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9496 6248 9548 6254
rect 9324 6174 9444 6202
rect 9496 6190 9548 6196
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 8956 4826 8984 5510
rect 9048 5234 9076 5646
rect 9140 5370 9168 6054
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4146 8432 4422
rect 8588 4282 8616 4762
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 6012 2514 6040 2790
rect 6656 2650 6684 2994
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6840 2446 6868 3062
rect 7300 2446 7328 3606
rect 7760 3466 7788 3878
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 3194 7604 3334
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7576 2446 7604 3130
rect 8496 2922 8524 4082
rect 8588 3126 8616 4218
rect 8864 4146 8892 4558
rect 9232 4486 9260 6054
rect 9416 5846 9444 6174
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5914 9536 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9416 5234 9444 5782
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9600 4486 9628 7890
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 6390 9720 7346
rect 9784 7290 9812 10560
rect 9876 10470 9904 10662
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10048 10668 10100 10674
rect 10100 10628 10180 10656
rect 10048 10610 10100 10616
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10062 9904 10406
rect 9968 10198 9996 10610
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9864 10056 9916 10062
rect 9956 10056 10008 10062
rect 9864 9998 9916 10004
rect 9954 10024 9956 10033
rect 10008 10024 10010 10033
rect 9876 8906 9904 9998
rect 9954 9959 10010 9968
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7478 9904 7822
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9784 7262 9904 7290
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6390 9812 7142
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9876 5914 9904 7262
rect 9968 6644 9996 9959
rect 10060 9586 10088 10474
rect 10152 10062 10180 10628
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10336 9722 10364 10746
rect 10428 10742 10456 11183
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10520 10606 10548 11319
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10612 10452 10640 11562
rect 11348 11558 11376 12406
rect 11532 12374 11560 12786
rect 11624 12782 11652 13126
rect 12084 12986 12112 13126
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11886 12880 11942 12889
rect 11886 12815 11942 12824
rect 12072 12844 12124 12850
rect 11900 12782 11928 12815
rect 12072 12786 12124 12792
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11624 12442 11652 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11610 12336 11666 12345
rect 11610 12271 11666 12280
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10784 11144 10836 11150
rect 10782 11112 10784 11121
rect 10968 11144 11020 11150
rect 10836 11112 10838 11121
rect 10782 11047 10838 11056
rect 10966 11112 10968 11121
rect 11060 11144 11112 11150
rect 11020 11112 11022 11121
rect 11060 11086 11112 11092
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 10966 11047 11022 11056
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10810 10732 10950
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10796 10674 10824 11047
rect 11072 11014 11100 11086
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10916 10908 11292 10917
rect 10972 10906 10996 10908
rect 11052 10906 11076 10908
rect 11132 10906 11156 10908
rect 11212 10906 11236 10908
rect 10972 10854 10982 10906
rect 11226 10854 11236 10906
rect 10972 10852 10996 10854
rect 11052 10852 11076 10854
rect 11132 10852 11156 10854
rect 11212 10852 11236 10854
rect 10916 10843 11292 10852
rect 11348 10810 11376 11086
rect 11440 11082 11468 12106
rect 11532 11898 11560 12174
rect 11624 11898 11652 12271
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11518 11792 11574 11801
rect 11716 11778 11744 12378
rect 11574 11750 11744 11778
rect 11518 11727 11574 11736
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11532 10810 11560 11727
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11624 10810 11652 11630
rect 11716 11558 11744 11630
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11808 11354 11836 12718
rect 11888 12368 11940 12374
rect 11886 12336 11888 12345
rect 11980 12368 12032 12374
rect 11940 12336 11942 12345
rect 11980 12310 12032 12316
rect 11886 12271 11942 12280
rect 11888 12232 11940 12238
rect 11886 12200 11888 12209
rect 11940 12200 11942 12209
rect 11886 12135 11942 12144
rect 11992 11762 12020 12310
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10704 10577 10732 10610
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10612 10424 10732 10452
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10060 8906 10088 9522
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 8090 10088 8842
rect 10152 8838 10180 9046
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10244 7546 10272 9522
rect 10336 9178 10364 9522
rect 10428 9178 10456 9522
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10336 7886 10364 8978
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10244 7002 10272 7142
rect 10336 7002 10364 7686
rect 10428 7342 10456 8774
rect 10520 8634 10548 9930
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 8838 10640 9862
rect 10704 9489 10732 10424
rect 10796 9994 10824 10610
rect 11256 10282 11284 10678
rect 11256 10254 11376 10282
rect 11348 10169 11376 10254
rect 11428 10192 11480 10198
rect 11334 10160 11390 10169
rect 11428 10134 11480 10140
rect 11334 10095 11390 10104
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10916 9820 11292 9829
rect 10972 9818 10996 9820
rect 11052 9818 11076 9820
rect 11132 9818 11156 9820
rect 11212 9818 11236 9820
rect 10972 9766 10982 9818
rect 11226 9766 11236 9818
rect 10972 9764 10996 9766
rect 11052 9764 11076 9766
rect 11132 9764 11156 9766
rect 11212 9764 11236 9766
rect 10916 9755 11292 9764
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10782 9616 10838 9625
rect 10782 9551 10838 9560
rect 10690 9480 10746 9489
rect 10690 9415 10746 9424
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9042 10732 9318
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10232 6792 10284 6798
rect 10152 6752 10232 6780
rect 10152 6644 10180 6752
rect 10232 6734 10284 6740
rect 9968 6616 10180 6644
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9692 4826 9720 5170
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9232 4146 9260 4422
rect 9692 4282 9720 4490
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9784 4146 9812 5510
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 8864 3466 8892 4082
rect 8956 3942 8984 4082
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8680 3194 8708 3402
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3194 8800 3334
rect 8956 3194 8984 3878
rect 9048 3466 9076 3878
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 9876 2446 9904 5510
rect 9968 4622 9996 6326
rect 10060 6186 10088 6616
rect 10336 6322 10364 6938
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10152 4622 10180 6190
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10336 5710 10364 5850
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10244 5370 10272 5646
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10336 5234 10364 5646
rect 10428 5234 10456 6054
rect 10520 5710 10548 8570
rect 10612 8090 10640 8774
rect 10796 8498 10824 9551
rect 10888 8974 10916 9658
rect 11348 9654 11376 10095
rect 11336 9648 11388 9654
rect 10966 9616 11022 9625
rect 11336 9590 11388 9596
rect 10966 9551 10968 9560
rect 11020 9551 11022 9560
rect 10968 9522 11020 9528
rect 10966 9480 11022 9489
rect 10966 9415 10968 9424
rect 11020 9415 11022 9424
rect 10968 9386 11020 9392
rect 10980 9178 11008 9386
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11072 8974 11100 9114
rect 11348 8974 11376 9590
rect 11440 8974 11468 10134
rect 11532 9518 11560 10746
rect 11900 10656 11928 10950
rect 11992 10810 12020 11698
rect 12084 11150 12112 12786
rect 12176 12714 12204 13212
rect 12256 13194 12308 13200
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12850 12388 13126
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12176 11762 12204 12650
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12268 12238 12296 12582
rect 12256 12232 12308 12238
rect 12440 12232 12492 12238
rect 12256 12174 12308 12180
rect 12360 12192 12440 12220
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11778 12296 12038
rect 12360 11898 12388 12192
rect 12440 12174 12492 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11898 12480 12038
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12164 11756 12216 11762
rect 12268 11750 12388 11778
rect 12164 11698 12216 11704
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11808 10628 11928 10656
rect 11978 10704 12034 10713
rect 12084 10674 12112 11086
rect 11978 10639 12034 10648
rect 12072 10668 12124 10674
rect 11808 10470 11836 10628
rect 11992 10606 12020 10639
rect 12072 10610 12124 10616
rect 11980 10600 12032 10606
rect 11900 10560 11980 10588
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 9926 11836 10406
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11532 9178 11560 9454
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 10916 8732 11292 8741
rect 10972 8730 10996 8732
rect 11052 8730 11076 8732
rect 11132 8730 11156 8732
rect 11212 8730 11236 8732
rect 10972 8678 10982 8730
rect 11226 8678 11236 8730
rect 10972 8676 10996 8678
rect 11052 8676 11076 8678
rect 11132 8676 11156 8678
rect 11212 8676 11236 8678
rect 10916 8667 11292 8676
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10796 7886 10824 8434
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10612 7410 10640 7754
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 10916 7644 11292 7653
rect 10972 7642 10996 7644
rect 11052 7642 11076 7644
rect 11132 7642 11156 7644
rect 11212 7642 11236 7644
rect 10972 7590 10982 7642
rect 11226 7590 11236 7642
rect 10972 7588 10996 7590
rect 11052 7588 11076 7590
rect 11132 7588 11156 7590
rect 11212 7588 11236 7590
rect 10916 7579 11292 7588
rect 11060 7540 11112 7546
rect 11348 7528 11376 7686
rect 11440 7546 11468 8910
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11060 7482 11112 7488
rect 11164 7500 11376 7528
rect 11428 7540 11480 7546
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 7002 10916 7142
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10612 6474 10640 6870
rect 10692 6792 10744 6798
rect 10690 6760 10692 6769
rect 10744 6760 10746 6769
rect 10690 6695 10746 6704
rect 10704 6644 10732 6695
rect 11072 6644 11100 7482
rect 11164 6934 11192 7500
rect 11428 7482 11480 7488
rect 11532 7410 11560 7890
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10704 6616 11100 6644
rect 10916 6556 11292 6565
rect 10972 6554 10996 6556
rect 11052 6554 11076 6556
rect 11132 6554 11156 6556
rect 11212 6554 11236 6556
rect 10972 6502 10982 6554
rect 11226 6502 11236 6554
rect 10972 6500 10996 6502
rect 11052 6500 11076 6502
rect 11132 6500 11156 6502
rect 11212 6500 11236 6502
rect 10916 6491 11292 6500
rect 10612 6446 10824 6474
rect 11348 6458 11376 7278
rect 11428 6928 11480 6934
rect 11532 6916 11560 7346
rect 11480 6888 11560 6916
rect 11428 6870 11480 6876
rect 11428 6786 11480 6792
rect 11428 6728 11480 6734
rect 10796 6338 10824 6446
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 10796 6322 11100 6338
rect 10600 6316 10652 6322
rect 10796 6316 11112 6322
rect 10796 6310 11060 6316
rect 10600 6258 10652 6264
rect 11440 6304 11468 6728
rect 11532 6322 11560 6888
rect 11060 6258 11112 6264
rect 11256 6276 11468 6304
rect 11520 6316 11572 6322
rect 10612 5846 10640 6258
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 11256 5574 11284 6276
rect 11520 6258 11572 6264
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10916 5468 11292 5477
rect 10972 5466 10996 5468
rect 11052 5466 11076 5468
rect 11132 5466 11156 5468
rect 11212 5466 11236 5468
rect 10972 5414 10982 5466
rect 11226 5414 11236 5466
rect 10972 5412 10996 5414
rect 11052 5412 11076 5414
rect 11132 5412 11156 5414
rect 11212 5412 11236 5414
rect 10916 5403 11292 5412
rect 11348 5234 11376 6054
rect 11440 5234 11468 6122
rect 11716 5846 11744 9318
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7002 11836 7822
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11900 6322 11928 10560
rect 11980 10542 12032 10548
rect 12084 9722 12112 10610
rect 12176 10266 12204 11698
rect 12360 11286 12388 11750
rect 12438 11384 12494 11393
rect 12438 11319 12440 11328
rect 12492 11319 12494 11328
rect 12440 11290 12492 11296
rect 12348 11280 12400 11286
rect 12544 11257 12572 12582
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12348 11222 12400 11228
rect 12530 11248 12586 11257
rect 12530 11183 12586 11192
rect 12544 11150 12572 11183
rect 12532 11144 12584 11150
rect 12346 11112 12402 11121
rect 12532 11086 12584 11092
rect 12346 11047 12402 11056
rect 12360 11014 12388 11047
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12176 9042 12204 10202
rect 12360 9382 12388 10950
rect 12544 10606 12572 10950
rect 12636 10810 12664 12174
rect 12728 12170 12756 12718
rect 13280 12345 13308 14214
rect 13266 12336 13322 12345
rect 13266 12271 13322 12280
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12728 10674 12756 12106
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9654 12480 10406
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12728 9450 12756 10610
rect 12820 10198 12848 12038
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13188 11354 13216 11494
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13556 11286 13584 11494
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12912 10606 12940 11086
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 8090 12020 8842
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 8498 13584 8774
rect 14200 8566 14228 16589
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12176 7954 12204 8230
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12452 7886 12480 8434
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12084 7410 12112 7822
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7410 12572 7686
rect 12820 7410 12848 7754
rect 12912 7410 12940 7890
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6798 12020 7142
rect 12084 6798 12112 7346
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12084 6118 12112 6734
rect 12820 6662 12848 7346
rect 12912 6798 12940 7346
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6254 12848 6598
rect 12912 6322 12940 6734
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 4758 10272 4966
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10336 4690 10364 5170
rect 10428 4826 10456 5170
rect 11532 5166 11560 5510
rect 12912 5370 12940 6258
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9968 4078 9996 4150
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10322 4040 10378 4049
rect 9968 3534 9996 4014
rect 10322 3975 10378 3984
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10336 3194 10364 3975
rect 10704 3534 10732 4422
rect 10916 4380 11292 4389
rect 10972 4378 10996 4380
rect 11052 4378 11076 4380
rect 11132 4378 11156 4380
rect 11212 4378 11236 4380
rect 10972 4326 10982 4378
rect 11226 4326 11236 4378
rect 10972 4324 10996 4326
rect 11052 4324 11076 4326
rect 11132 4324 11156 4326
rect 11212 4324 11236 4326
rect 10916 4315 11292 4324
rect 11348 3942 11376 4966
rect 11532 4690 11560 5102
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4214 11560 4626
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11808 3738 11836 4558
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13464 4282 13492 4490
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10916 3292 11292 3301
rect 10972 3290 10996 3292
rect 11052 3290 11076 3292
rect 11132 3290 11156 3292
rect 11212 3290 11236 3292
rect 10972 3238 10982 3290
rect 11226 3238 11236 3290
rect 10972 3236 10996 3238
rect 11052 3236 11076 3238
rect 11132 3236 11156 3238
rect 11212 3236 11236 3238
rect 10916 3227 11292 3236
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10428 2446 10456 2790
rect 12084 2446 12112 3878
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12176 2446 12204 3674
rect 13556 2650 13584 4082
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 1032 2304 1084 2310
rect 2320 2304 2372 2310
rect 1032 2246 1084 2252
rect 2240 2264 2320 2292
rect 1044 800 1072 2246
rect 2240 800 2268 2264
rect 2320 2246 2372 2252
rect 3424 2304 3476 2310
rect 4712 2304 4764 2310
rect 3424 2246 3476 2252
rect 4632 2264 4712 2292
rect 3436 800 3464 2246
rect 4632 800 4660 2264
rect 5908 2304 5960 2310
rect 4712 2246 4764 2252
rect 5828 2264 5908 2292
rect 4916 2204 5292 2213
rect 4972 2202 4996 2204
rect 5052 2202 5076 2204
rect 5132 2202 5156 2204
rect 5212 2202 5236 2204
rect 4972 2150 4982 2202
rect 5226 2150 5236 2202
rect 4972 2148 4996 2150
rect 5052 2148 5076 2150
rect 5132 2148 5156 2150
rect 5212 2148 5236 2150
rect 4916 2139 5292 2148
rect 5828 800 5856 2264
rect 5908 2246 5960 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 7116 1170 7144 2246
rect 7024 1142 7144 1170
rect 7024 800 7052 1142
rect 8220 800 8248 2246
rect 9508 1170 9536 2246
rect 10704 1170 10732 2246
rect 10916 2204 11292 2213
rect 10972 2202 10996 2204
rect 11052 2202 11076 2204
rect 11132 2202 11156 2204
rect 11212 2202 11236 2204
rect 10972 2150 10982 2202
rect 11226 2150 11236 2202
rect 10972 2148 10996 2150
rect 11052 2148 11076 2150
rect 11132 2148 11156 2150
rect 11212 2148 11236 2150
rect 10916 2139 11292 2148
rect 11900 1170 11928 2246
rect 13096 1170 13124 2246
rect 9416 1142 9536 1170
rect 10612 1142 10732 1170
rect 11808 1142 11928 1170
rect 13004 1142 13124 1170
rect 9416 800 9444 1142
rect 10612 800 10640 1142
rect 11808 800 11836 1142
rect 13004 800 13032 1142
rect 14200 800 14228 2382
rect 1030 0 1086 800
rect 2226 0 2282 800
rect 3422 0 3478 800
rect 4618 0 4674 800
rect 5814 0 5870 800
rect 7010 0 7066 800
rect 8206 0 8262 800
rect 9402 0 9458 800
rect 10598 0 10654 800
rect 11794 0 11850 800
rect 12990 0 13046 800
rect 14186 0 14242 800
<< via2 >>
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 3422 11192 3478 11248
rect 3238 11056 3294 11112
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 2318 9016 2374 9072
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 4250 12180 4252 12200
rect 4252 12180 4304 12200
rect 4304 12180 4306 12200
rect 4250 12144 4306 12180
rect 3606 9560 3662 9616
rect 3790 10104 3846 10160
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 3238 5480 3294 5536
rect 4916 14170 4972 14172
rect 4996 14170 5052 14172
rect 5076 14170 5132 14172
rect 5156 14170 5212 14172
rect 5236 14170 5292 14172
rect 4916 14118 4918 14170
rect 4918 14118 4970 14170
rect 4970 14118 4972 14170
rect 4996 14118 5034 14170
rect 5034 14118 5046 14170
rect 5046 14118 5052 14170
rect 5076 14118 5098 14170
rect 5098 14118 5110 14170
rect 5110 14118 5132 14170
rect 5156 14118 5162 14170
rect 5162 14118 5174 14170
rect 5174 14118 5212 14170
rect 5236 14118 5238 14170
rect 5238 14118 5290 14170
rect 5290 14118 5292 14170
rect 4916 14116 4972 14118
rect 4996 14116 5052 14118
rect 5076 14116 5132 14118
rect 5156 14116 5212 14118
rect 5236 14116 5292 14118
rect 4916 13082 4972 13084
rect 4996 13082 5052 13084
rect 5076 13082 5132 13084
rect 5156 13082 5212 13084
rect 5236 13082 5292 13084
rect 4916 13030 4918 13082
rect 4918 13030 4970 13082
rect 4970 13030 4972 13082
rect 4996 13030 5034 13082
rect 5034 13030 5046 13082
rect 5046 13030 5052 13082
rect 5076 13030 5098 13082
rect 5098 13030 5110 13082
rect 5110 13030 5132 13082
rect 5156 13030 5162 13082
rect 5162 13030 5174 13082
rect 5174 13030 5212 13082
rect 5236 13030 5238 13082
rect 5238 13030 5290 13082
rect 5290 13030 5292 13082
rect 4916 13028 4972 13030
rect 4996 13028 5052 13030
rect 5076 13028 5132 13030
rect 5156 13028 5212 13030
rect 5236 13028 5292 13030
rect 4916 11994 4972 11996
rect 4996 11994 5052 11996
rect 5076 11994 5132 11996
rect 5156 11994 5212 11996
rect 5236 11994 5292 11996
rect 4916 11942 4918 11994
rect 4918 11942 4970 11994
rect 4970 11942 4972 11994
rect 4996 11942 5034 11994
rect 5034 11942 5046 11994
rect 5046 11942 5052 11994
rect 5076 11942 5098 11994
rect 5098 11942 5110 11994
rect 5110 11942 5132 11994
rect 5156 11942 5162 11994
rect 5162 11942 5174 11994
rect 5174 11942 5212 11994
rect 5236 11942 5238 11994
rect 5238 11942 5290 11994
rect 5290 11942 5292 11994
rect 4916 11940 4972 11942
rect 4996 11940 5052 11942
rect 5076 11940 5132 11942
rect 5156 11940 5212 11942
rect 5236 11940 5292 11942
rect 4916 10906 4972 10908
rect 4996 10906 5052 10908
rect 5076 10906 5132 10908
rect 5156 10906 5212 10908
rect 5236 10906 5292 10908
rect 4916 10854 4918 10906
rect 4918 10854 4970 10906
rect 4970 10854 4972 10906
rect 4996 10854 5034 10906
rect 5034 10854 5046 10906
rect 5046 10854 5052 10906
rect 5076 10854 5098 10906
rect 5098 10854 5110 10906
rect 5110 10854 5132 10906
rect 5156 10854 5162 10906
rect 5162 10854 5174 10906
rect 5174 10854 5212 10906
rect 5236 10854 5238 10906
rect 5238 10854 5290 10906
rect 5290 10854 5292 10906
rect 4916 10852 4972 10854
rect 4996 10852 5052 10854
rect 5076 10852 5132 10854
rect 5156 10852 5212 10854
rect 5236 10852 5292 10854
rect 4618 9424 4674 9480
rect 3054 3984 3110 4040
rect 5262 9968 5318 10024
rect 4916 9818 4972 9820
rect 4996 9818 5052 9820
rect 5076 9818 5132 9820
rect 5156 9818 5212 9820
rect 5236 9818 5292 9820
rect 4916 9766 4918 9818
rect 4918 9766 4970 9818
rect 4970 9766 4972 9818
rect 4996 9766 5034 9818
rect 5034 9766 5046 9818
rect 5046 9766 5052 9818
rect 5076 9766 5098 9818
rect 5098 9766 5110 9818
rect 5110 9766 5132 9818
rect 5156 9766 5162 9818
rect 5162 9766 5174 9818
rect 5174 9766 5212 9818
rect 5236 9766 5238 9818
rect 5238 9766 5290 9818
rect 5290 9766 5292 9818
rect 4916 9764 4972 9766
rect 4996 9764 5052 9766
rect 5076 9764 5132 9766
rect 5156 9764 5212 9766
rect 5236 9764 5292 9766
rect 4894 9596 4896 9616
rect 4896 9596 4948 9616
rect 4948 9596 4950 9616
rect 4894 9560 4950 9596
rect 5078 9016 5134 9072
rect 5630 10548 5632 10568
rect 5632 10548 5684 10568
rect 5684 10548 5686 10568
rect 5630 10512 5686 10548
rect 4986 8880 5042 8936
rect 4916 8730 4972 8732
rect 4996 8730 5052 8732
rect 5076 8730 5132 8732
rect 5156 8730 5212 8732
rect 5236 8730 5292 8732
rect 4916 8678 4918 8730
rect 4918 8678 4970 8730
rect 4970 8678 4972 8730
rect 4996 8678 5034 8730
rect 5034 8678 5046 8730
rect 5046 8678 5052 8730
rect 5076 8678 5098 8730
rect 5098 8678 5110 8730
rect 5110 8678 5132 8730
rect 5156 8678 5162 8730
rect 5162 8678 5174 8730
rect 5174 8678 5212 8730
rect 5236 8678 5238 8730
rect 5238 8678 5290 8730
rect 5290 8678 5292 8730
rect 4916 8676 4972 8678
rect 4996 8676 5052 8678
rect 5076 8676 5132 8678
rect 5156 8676 5212 8678
rect 5236 8676 5292 8678
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 4916 7642 4972 7644
rect 4996 7642 5052 7644
rect 5076 7642 5132 7644
rect 5156 7642 5212 7644
rect 5236 7642 5292 7644
rect 4916 7590 4918 7642
rect 4918 7590 4970 7642
rect 4970 7590 4972 7642
rect 4996 7590 5034 7642
rect 5034 7590 5046 7642
rect 5046 7590 5052 7642
rect 5076 7590 5098 7642
rect 5098 7590 5110 7642
rect 5110 7590 5132 7642
rect 5156 7590 5162 7642
rect 5162 7590 5174 7642
rect 5174 7590 5212 7642
rect 5236 7590 5238 7642
rect 5238 7590 5290 7642
rect 5290 7590 5292 7642
rect 4916 7588 4972 7590
rect 4996 7588 5052 7590
rect 5076 7588 5132 7590
rect 5156 7588 5212 7590
rect 5236 7588 5292 7590
rect 4916 6554 4972 6556
rect 4996 6554 5052 6556
rect 5076 6554 5132 6556
rect 5156 6554 5212 6556
rect 5236 6554 5292 6556
rect 4916 6502 4918 6554
rect 4918 6502 4970 6554
rect 4970 6502 4972 6554
rect 4996 6502 5034 6554
rect 5034 6502 5046 6554
rect 5046 6502 5052 6554
rect 5076 6502 5098 6554
rect 5098 6502 5110 6554
rect 5110 6502 5132 6554
rect 5156 6502 5162 6554
rect 5162 6502 5174 6554
rect 5174 6502 5212 6554
rect 5236 6502 5238 6554
rect 5238 6502 5290 6554
rect 5290 6502 5292 6554
rect 4916 6500 4972 6502
rect 4996 6500 5052 6502
rect 5076 6500 5132 6502
rect 5156 6500 5212 6502
rect 5236 6500 5292 6502
rect 4916 5466 4972 5468
rect 4996 5466 5052 5468
rect 5076 5466 5132 5468
rect 5156 5466 5212 5468
rect 5236 5466 5292 5468
rect 4916 5414 4918 5466
rect 4918 5414 4970 5466
rect 4970 5414 4972 5466
rect 4996 5414 5034 5466
rect 5034 5414 5046 5466
rect 5046 5414 5052 5466
rect 5076 5414 5098 5466
rect 5098 5414 5110 5466
rect 5110 5414 5132 5466
rect 5156 5414 5162 5466
rect 5162 5414 5174 5466
rect 5174 5414 5212 5466
rect 5236 5414 5238 5466
rect 5238 5414 5290 5466
rect 5290 5414 5292 5466
rect 4916 5412 4972 5414
rect 4996 5412 5052 5414
rect 5076 5412 5132 5414
rect 5156 5412 5212 5414
rect 5236 5412 5292 5414
rect 4916 4378 4972 4380
rect 4996 4378 5052 4380
rect 5076 4378 5132 4380
rect 5156 4378 5212 4380
rect 5236 4378 5292 4380
rect 4916 4326 4918 4378
rect 4918 4326 4970 4378
rect 4970 4326 4972 4378
rect 4996 4326 5034 4378
rect 5034 4326 5046 4378
rect 5046 4326 5052 4378
rect 5076 4326 5098 4378
rect 5098 4326 5110 4378
rect 5110 4326 5132 4378
rect 5156 4326 5162 4378
rect 5162 4326 5174 4378
rect 5174 4326 5212 4378
rect 5236 4326 5238 4378
rect 5238 4326 5290 4378
rect 5290 4326 5292 4378
rect 4916 4324 4972 4326
rect 4996 4324 5052 4326
rect 5076 4324 5132 4326
rect 5156 4324 5212 4326
rect 5236 4324 5292 4326
rect 7378 10648 7434 10704
rect 6826 9444 6882 9480
rect 6826 9424 6828 9444
rect 6828 9424 6880 9444
rect 6880 9424 6882 9444
rect 6734 9016 6790 9072
rect 7194 9696 7250 9752
rect 7010 9596 7012 9616
rect 7012 9596 7064 9616
rect 7064 9596 7066 9616
rect 7010 9560 7066 9596
rect 7102 8900 7158 8936
rect 7102 8880 7104 8900
rect 7104 8880 7156 8900
rect 7156 8880 7158 8900
rect 7010 6196 7012 6216
rect 7012 6196 7064 6216
rect 7064 6196 7066 6216
rect 7010 6160 7066 6196
rect 4916 3290 4972 3292
rect 4996 3290 5052 3292
rect 5076 3290 5132 3292
rect 5156 3290 5212 3292
rect 5236 3290 5292 3292
rect 4916 3238 4918 3290
rect 4918 3238 4970 3290
rect 4970 3238 4972 3290
rect 4996 3238 5034 3290
rect 5034 3238 5046 3290
rect 5046 3238 5052 3290
rect 5076 3238 5098 3290
rect 5098 3238 5110 3290
rect 5110 3238 5132 3290
rect 5156 3238 5162 3290
rect 5162 3238 5174 3290
rect 5174 3238 5212 3290
rect 5236 3238 5238 3290
rect 5238 3238 5290 3290
rect 5290 3238 5292 3290
rect 4916 3236 4972 3238
rect 4996 3236 5052 3238
rect 5076 3236 5132 3238
rect 5156 3236 5212 3238
rect 5236 3236 5292 3238
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 10916 14170 10972 14172
rect 10996 14170 11052 14172
rect 11076 14170 11132 14172
rect 11156 14170 11212 14172
rect 11236 14170 11292 14172
rect 10916 14118 10918 14170
rect 10918 14118 10970 14170
rect 10970 14118 10972 14170
rect 10996 14118 11034 14170
rect 11034 14118 11046 14170
rect 11046 14118 11052 14170
rect 11076 14118 11098 14170
rect 11098 14118 11110 14170
rect 11110 14118 11132 14170
rect 11156 14118 11162 14170
rect 11162 14118 11174 14170
rect 11174 14118 11212 14170
rect 11236 14118 11238 14170
rect 11238 14118 11290 14170
rect 11290 14118 11292 14170
rect 10916 14116 10972 14118
rect 10996 14116 11052 14118
rect 11076 14116 11132 14118
rect 11156 14116 11212 14118
rect 11236 14116 11292 14118
rect 11518 13776 11574 13832
rect 12254 13776 12310 13832
rect 10138 13640 10194 13696
rect 9862 12860 9864 12880
rect 9864 12860 9916 12880
rect 9916 12860 9918 12880
rect 9126 12280 9182 12336
rect 9862 12824 9918 12860
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 7838 10668 7894 10704
rect 7838 10648 7840 10668
rect 7840 10648 7892 10668
rect 7892 10648 7894 10668
rect 8114 10548 8116 10568
rect 8116 10548 8168 10568
rect 8168 10548 8170 10568
rect 8114 10512 8170 10548
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 8298 10104 8354 10160
rect 8390 9868 8392 9888
rect 8392 9868 8444 9888
rect 8444 9868 8446 9888
rect 8390 9832 8446 9868
rect 8206 9696 8262 9752
rect 8114 9460 8116 9480
rect 8116 9460 8168 9480
rect 8168 9460 8170 9480
rect 8114 9424 8170 9460
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 8666 9596 8668 9616
rect 8668 9596 8720 9616
rect 8720 9596 8722 9616
rect 8666 9560 8722 9596
rect 8758 9460 8760 9480
rect 8760 9460 8812 9480
rect 8812 9460 8814 9480
rect 8758 9424 8814 9460
rect 10916 13082 10972 13084
rect 10996 13082 11052 13084
rect 11076 13082 11132 13084
rect 11156 13082 11212 13084
rect 11236 13082 11292 13084
rect 10916 13030 10918 13082
rect 10918 13030 10970 13082
rect 10970 13030 10972 13082
rect 10996 13030 11034 13082
rect 11034 13030 11046 13082
rect 11046 13030 11052 13082
rect 11076 13030 11098 13082
rect 11098 13030 11110 13082
rect 11110 13030 11132 13082
rect 11156 13030 11162 13082
rect 11162 13030 11174 13082
rect 11174 13030 11212 13082
rect 11236 13030 11238 13082
rect 11238 13030 11290 13082
rect 11290 13030 11292 13082
rect 10916 13028 10972 13030
rect 10996 13028 11052 13030
rect 11076 13028 11132 13030
rect 11156 13028 11212 13030
rect 11236 13028 11292 13030
rect 9770 11756 9826 11792
rect 9770 11736 9772 11756
rect 9772 11736 9824 11756
rect 9824 11736 9826 11756
rect 9954 11056 10010 11112
rect 11242 12316 11244 12336
rect 11244 12316 11296 12336
rect 11296 12316 11298 12336
rect 11242 12280 11298 12316
rect 10916 11994 10972 11996
rect 10996 11994 11052 11996
rect 11076 11994 11132 11996
rect 11156 11994 11212 11996
rect 11236 11994 11292 11996
rect 10916 11942 10918 11994
rect 10918 11942 10970 11994
rect 10970 11942 10972 11994
rect 10996 11942 11034 11994
rect 11034 11942 11046 11994
rect 11046 11942 11052 11994
rect 11076 11942 11098 11994
rect 11098 11942 11110 11994
rect 11110 11942 11132 11994
rect 11156 11942 11162 11994
rect 11162 11942 11174 11994
rect 11174 11942 11212 11994
rect 11236 11942 11238 11994
rect 11238 11942 11290 11994
rect 11290 11942 11292 11994
rect 10916 11940 10972 11942
rect 10996 11940 11052 11942
rect 11076 11940 11132 11942
rect 11156 11940 11212 11942
rect 11236 11940 11292 11942
rect 10506 11328 10562 11384
rect 10414 11192 10470 11248
rect 9310 9832 9366 9888
rect 8574 9016 8630 9072
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 8206 6704 8262 6760
rect 8482 6976 8538 7032
rect 9402 6996 9458 7032
rect 9402 6976 9404 6996
rect 9404 6976 9456 6996
rect 9456 6976 9458 6996
rect 7746 6180 7802 6216
rect 7746 6160 7748 6180
rect 7748 6160 7800 6180
rect 7800 6160 7802 6180
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 9954 10004 9956 10024
rect 9956 10004 10008 10024
rect 10008 10004 10010 10024
rect 9954 9968 10010 10004
rect 11886 12824 11942 12880
rect 11610 12280 11666 12336
rect 10782 11092 10784 11112
rect 10784 11092 10836 11112
rect 10836 11092 10838 11112
rect 10782 11056 10838 11092
rect 10966 11092 10968 11112
rect 10968 11092 11020 11112
rect 11020 11092 11022 11112
rect 10966 11056 11022 11092
rect 10916 10906 10972 10908
rect 10996 10906 11052 10908
rect 11076 10906 11132 10908
rect 11156 10906 11212 10908
rect 11236 10906 11292 10908
rect 10916 10854 10918 10906
rect 10918 10854 10970 10906
rect 10970 10854 10972 10906
rect 10996 10854 11034 10906
rect 11034 10854 11046 10906
rect 11046 10854 11052 10906
rect 11076 10854 11098 10906
rect 11098 10854 11110 10906
rect 11110 10854 11132 10906
rect 11156 10854 11162 10906
rect 11162 10854 11174 10906
rect 11174 10854 11212 10906
rect 11236 10854 11238 10906
rect 11238 10854 11290 10906
rect 11290 10854 11292 10906
rect 10916 10852 10972 10854
rect 10996 10852 11052 10854
rect 11076 10852 11132 10854
rect 11156 10852 11212 10854
rect 11236 10852 11292 10854
rect 11518 11736 11574 11792
rect 11886 12316 11888 12336
rect 11888 12316 11940 12336
rect 11940 12316 11942 12336
rect 11886 12280 11942 12316
rect 11886 12180 11888 12200
rect 11888 12180 11940 12200
rect 11940 12180 11942 12200
rect 11886 12144 11942 12180
rect 10690 10512 10746 10568
rect 11334 10104 11390 10160
rect 10916 9818 10972 9820
rect 10996 9818 11052 9820
rect 11076 9818 11132 9820
rect 11156 9818 11212 9820
rect 11236 9818 11292 9820
rect 10916 9766 10918 9818
rect 10918 9766 10970 9818
rect 10970 9766 10972 9818
rect 10996 9766 11034 9818
rect 11034 9766 11046 9818
rect 11046 9766 11052 9818
rect 11076 9766 11098 9818
rect 11098 9766 11110 9818
rect 11110 9766 11132 9818
rect 11156 9766 11162 9818
rect 11162 9766 11174 9818
rect 11174 9766 11212 9818
rect 11236 9766 11238 9818
rect 11238 9766 11290 9818
rect 11290 9766 11292 9818
rect 10916 9764 10972 9766
rect 10996 9764 11052 9766
rect 11076 9764 11132 9766
rect 11156 9764 11212 9766
rect 11236 9764 11292 9766
rect 10782 9560 10838 9616
rect 10690 9424 10746 9480
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 10966 9580 11022 9616
rect 10966 9560 10968 9580
rect 10968 9560 11020 9580
rect 11020 9560 11022 9580
rect 10966 9444 11022 9480
rect 10966 9424 10968 9444
rect 10968 9424 11020 9444
rect 11020 9424 11022 9444
rect 11978 10648 12034 10704
rect 10916 8730 10972 8732
rect 10996 8730 11052 8732
rect 11076 8730 11132 8732
rect 11156 8730 11212 8732
rect 11236 8730 11292 8732
rect 10916 8678 10918 8730
rect 10918 8678 10970 8730
rect 10970 8678 10972 8730
rect 10996 8678 11034 8730
rect 11034 8678 11046 8730
rect 11046 8678 11052 8730
rect 11076 8678 11098 8730
rect 11098 8678 11110 8730
rect 11110 8678 11132 8730
rect 11156 8678 11162 8730
rect 11162 8678 11174 8730
rect 11174 8678 11212 8730
rect 11236 8678 11238 8730
rect 11238 8678 11290 8730
rect 11290 8678 11292 8730
rect 10916 8676 10972 8678
rect 10996 8676 11052 8678
rect 11076 8676 11132 8678
rect 11156 8676 11212 8678
rect 11236 8676 11292 8678
rect 10916 7642 10972 7644
rect 10996 7642 11052 7644
rect 11076 7642 11132 7644
rect 11156 7642 11212 7644
rect 11236 7642 11292 7644
rect 10916 7590 10918 7642
rect 10918 7590 10970 7642
rect 10970 7590 10972 7642
rect 10996 7590 11034 7642
rect 11034 7590 11046 7642
rect 11046 7590 11052 7642
rect 11076 7590 11098 7642
rect 11098 7590 11110 7642
rect 11110 7590 11132 7642
rect 11156 7590 11162 7642
rect 11162 7590 11174 7642
rect 11174 7590 11212 7642
rect 11236 7590 11238 7642
rect 11238 7590 11290 7642
rect 11290 7590 11292 7642
rect 10916 7588 10972 7590
rect 10996 7588 11052 7590
rect 11076 7588 11132 7590
rect 11156 7588 11212 7590
rect 11236 7588 11292 7590
rect 10690 6740 10692 6760
rect 10692 6740 10744 6760
rect 10744 6740 10746 6760
rect 10690 6704 10746 6740
rect 10916 6554 10972 6556
rect 10996 6554 11052 6556
rect 11076 6554 11132 6556
rect 11156 6554 11212 6556
rect 11236 6554 11292 6556
rect 10916 6502 10918 6554
rect 10918 6502 10970 6554
rect 10970 6502 10972 6554
rect 10996 6502 11034 6554
rect 11034 6502 11046 6554
rect 11046 6502 11052 6554
rect 11076 6502 11098 6554
rect 11098 6502 11110 6554
rect 11110 6502 11132 6554
rect 11156 6502 11162 6554
rect 11162 6502 11174 6554
rect 11174 6502 11212 6554
rect 11236 6502 11238 6554
rect 11238 6502 11290 6554
rect 11290 6502 11292 6554
rect 10916 6500 10972 6502
rect 10996 6500 11052 6502
rect 11076 6500 11132 6502
rect 11156 6500 11212 6502
rect 11236 6500 11292 6502
rect 10916 5466 10972 5468
rect 10996 5466 11052 5468
rect 11076 5466 11132 5468
rect 11156 5466 11212 5468
rect 11236 5466 11292 5468
rect 10916 5414 10918 5466
rect 10918 5414 10970 5466
rect 10970 5414 10972 5466
rect 10996 5414 11034 5466
rect 11034 5414 11046 5466
rect 11046 5414 11052 5466
rect 11076 5414 11098 5466
rect 11098 5414 11110 5466
rect 11110 5414 11132 5466
rect 11156 5414 11162 5466
rect 11162 5414 11174 5466
rect 11174 5414 11212 5466
rect 11236 5414 11238 5466
rect 11238 5414 11290 5466
rect 11290 5414 11292 5466
rect 10916 5412 10972 5414
rect 10996 5412 11052 5414
rect 11076 5412 11132 5414
rect 11156 5412 11212 5414
rect 11236 5412 11292 5414
rect 12438 11348 12494 11384
rect 12438 11328 12440 11348
rect 12440 11328 12492 11348
rect 12492 11328 12494 11348
rect 12530 11192 12586 11248
rect 12346 11056 12402 11112
rect 13266 12280 13322 12336
rect 10322 3984 10378 4040
rect 10916 4378 10972 4380
rect 10996 4378 11052 4380
rect 11076 4378 11132 4380
rect 11156 4378 11212 4380
rect 11236 4378 11292 4380
rect 10916 4326 10918 4378
rect 10918 4326 10970 4378
rect 10970 4326 10972 4378
rect 10996 4326 11034 4378
rect 11034 4326 11046 4378
rect 11046 4326 11052 4378
rect 11076 4326 11098 4378
rect 11098 4326 11110 4378
rect 11110 4326 11132 4378
rect 11156 4326 11162 4378
rect 11162 4326 11174 4378
rect 11174 4326 11212 4378
rect 11236 4326 11238 4378
rect 11238 4326 11290 4378
rect 11290 4326 11292 4378
rect 10916 4324 10972 4326
rect 10996 4324 11052 4326
rect 11076 4324 11132 4326
rect 11156 4324 11212 4326
rect 11236 4324 11292 4326
rect 10916 3290 10972 3292
rect 10996 3290 11052 3292
rect 11076 3290 11132 3292
rect 11156 3290 11212 3292
rect 11236 3290 11292 3292
rect 10916 3238 10918 3290
rect 10918 3238 10970 3290
rect 10970 3238 10972 3290
rect 10996 3238 11034 3290
rect 11034 3238 11046 3290
rect 11046 3238 11052 3290
rect 11076 3238 11098 3290
rect 11098 3238 11110 3290
rect 11110 3238 11132 3290
rect 11156 3238 11162 3290
rect 11162 3238 11174 3290
rect 11174 3238 11212 3290
rect 11236 3238 11238 3290
rect 11238 3238 11290 3290
rect 11290 3238 11292 3290
rect 10916 3236 10972 3238
rect 10996 3236 11052 3238
rect 11076 3236 11132 3238
rect 11156 3236 11212 3238
rect 11236 3236 11292 3238
rect 4916 2202 4972 2204
rect 4996 2202 5052 2204
rect 5076 2202 5132 2204
rect 5156 2202 5212 2204
rect 5236 2202 5292 2204
rect 4916 2150 4918 2202
rect 4918 2150 4970 2202
rect 4970 2150 4972 2202
rect 4996 2150 5034 2202
rect 5034 2150 5046 2202
rect 5046 2150 5052 2202
rect 5076 2150 5098 2202
rect 5098 2150 5110 2202
rect 5110 2150 5132 2202
rect 5156 2150 5162 2202
rect 5162 2150 5174 2202
rect 5174 2150 5212 2202
rect 5236 2150 5238 2202
rect 5238 2150 5290 2202
rect 5290 2150 5292 2202
rect 4916 2148 4972 2150
rect 4996 2148 5052 2150
rect 5076 2148 5132 2150
rect 5156 2148 5212 2150
rect 5236 2148 5292 2150
rect 10916 2202 10972 2204
rect 10996 2202 11052 2204
rect 11076 2202 11132 2204
rect 11156 2202 11212 2204
rect 11236 2202 11292 2204
rect 10916 2150 10918 2202
rect 10918 2150 10970 2202
rect 10970 2150 10972 2202
rect 10996 2150 11034 2202
rect 11034 2150 11046 2202
rect 11046 2150 11052 2202
rect 11076 2150 11098 2202
rect 11098 2150 11110 2202
rect 11110 2150 11132 2202
rect 11156 2150 11162 2202
rect 11162 2150 11174 2202
rect 11174 2150 11212 2202
rect 11236 2150 11238 2202
rect 11238 2150 11290 2202
rect 11290 2150 11292 2202
rect 10916 2148 10972 2150
rect 10996 2148 11052 2150
rect 11076 2148 11132 2150
rect 11156 2148 11212 2150
rect 11236 2148 11292 2150
<< metal3 >>
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 4906 14176 5302 14177
rect 4906 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5302 14176
rect 4906 14111 5302 14112
rect 10906 14176 11302 14177
rect 10906 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11302 14176
rect 10906 14111 11302 14112
rect 10726 13772 10732 13836
rect 10796 13834 10802 13836
rect 11513 13834 11579 13837
rect 12249 13836 12315 13837
rect 12198 13834 12204 13836
rect 10796 13832 11579 13834
rect 10796 13776 11518 13832
rect 11574 13776 11579 13832
rect 10796 13774 11579 13776
rect 12158 13774 12204 13834
rect 12268 13832 12315 13836
rect 12310 13776 12315 13832
rect 10796 13772 10802 13774
rect 11513 13771 11579 13774
rect 12198 13772 12204 13774
rect 12268 13772 12315 13776
rect 12249 13771 12315 13772
rect 10133 13698 10199 13701
rect 10358 13698 10364 13700
rect 10133 13696 10364 13698
rect 10133 13640 10138 13696
rect 10194 13640 10364 13696
rect 10133 13638 10364 13640
rect 10133 13635 10199 13638
rect 10358 13636 10364 13638
rect 10428 13636 10434 13700
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 4906 13088 5302 13089
rect 4906 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5302 13088
rect 4906 13023 5302 13024
rect 10906 13088 11302 13089
rect 10906 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11302 13088
rect 10906 13023 11302 13024
rect 9857 12882 9923 12885
rect 11881 12882 11947 12885
rect 9857 12880 11947 12882
rect 9857 12824 9862 12880
rect 9918 12824 11886 12880
rect 11942 12824 11947 12880
rect 9857 12822 11947 12824
rect 9857 12819 9923 12822
rect 11881 12819 11947 12822
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 9121 12338 9187 12341
rect 11237 12338 11303 12341
rect 9121 12336 11303 12338
rect 9121 12280 9126 12336
rect 9182 12280 11242 12336
rect 11298 12280 11303 12336
rect 9121 12278 11303 12280
rect 9121 12275 9187 12278
rect 11237 12275 11303 12278
rect 11605 12338 11671 12341
rect 11881 12338 11947 12341
rect 13261 12338 13327 12341
rect 11605 12336 11947 12338
rect 11605 12280 11610 12336
rect 11666 12280 11886 12336
rect 11942 12280 11947 12336
rect 11605 12278 11947 12280
rect 11605 12275 11671 12278
rect 11881 12275 11947 12278
rect 12390 12336 13327 12338
rect 12390 12280 13266 12336
rect 13322 12280 13327 12336
rect 12390 12278 13327 12280
rect 4245 12202 4311 12205
rect 11881 12202 11947 12205
rect 12390 12202 12450 12278
rect 13261 12275 13327 12278
rect 4245 12200 12450 12202
rect 4245 12144 4250 12200
rect 4306 12144 11886 12200
rect 11942 12144 12450 12200
rect 4245 12142 12450 12144
rect 4245 12139 4311 12142
rect 11881 12139 11947 12142
rect 4906 12000 5302 12001
rect 4906 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5302 12000
rect 4906 11935 5302 11936
rect 10906 12000 11302 12001
rect 10906 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11302 12000
rect 10906 11935 11302 11936
rect 9765 11794 9831 11797
rect 11513 11794 11579 11797
rect 9765 11792 11579 11794
rect 9765 11736 9770 11792
rect 9826 11736 11518 11792
rect 11574 11736 11579 11792
rect 9765 11734 11579 11736
rect 9765 11731 9831 11734
rect 11513 11731 11579 11734
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 10501 11386 10567 11389
rect 12433 11386 12499 11389
rect 10501 11384 12499 11386
rect 10501 11328 10506 11384
rect 10562 11328 12438 11384
rect 12494 11328 12499 11384
rect 10501 11326 12499 11328
rect 10501 11323 10567 11326
rect 12433 11323 12499 11326
rect 3417 11252 3483 11253
rect 3366 11188 3372 11252
rect 3436 11250 3483 11252
rect 10409 11250 10475 11253
rect 12525 11250 12591 11253
rect 3436 11248 3528 11250
rect 3478 11192 3528 11248
rect 3436 11190 3528 11192
rect 10409 11248 12591 11250
rect 10409 11192 10414 11248
rect 10470 11192 12530 11248
rect 12586 11192 12591 11248
rect 10409 11190 12591 11192
rect 3436 11188 3483 11190
rect 3417 11187 3483 11188
rect 10409 11187 10475 11190
rect 12525 11187 12591 11190
rect 3233 11116 3299 11117
rect 3182 11052 3188 11116
rect 3252 11114 3299 11116
rect 9949 11114 10015 11117
rect 10777 11114 10843 11117
rect 3252 11112 3344 11114
rect 3294 11056 3344 11112
rect 3252 11054 3344 11056
rect 9949 11112 10843 11114
rect 9949 11056 9954 11112
rect 10010 11056 10782 11112
rect 10838 11056 10843 11112
rect 9949 11054 10843 11056
rect 3252 11052 3299 11054
rect 3233 11051 3299 11052
rect 9949 11051 10015 11054
rect 10777 11051 10843 11054
rect 10961 11114 11027 11117
rect 12341 11114 12407 11117
rect 10961 11112 12407 11114
rect 10961 11056 10966 11112
rect 11022 11056 12346 11112
rect 12402 11056 12407 11112
rect 10961 11054 12407 11056
rect 10961 11051 11027 11054
rect 12341 11051 12407 11054
rect 4906 10912 5302 10913
rect 4906 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5302 10912
rect 4906 10847 5302 10848
rect 10906 10912 11302 10913
rect 10906 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11302 10912
rect 10906 10847 11302 10848
rect 7373 10706 7439 10709
rect 7833 10706 7899 10709
rect 7373 10704 7899 10706
rect 7373 10648 7378 10704
rect 7434 10648 7838 10704
rect 7894 10648 7899 10704
rect 7373 10646 7899 10648
rect 7373 10643 7439 10646
rect 7833 10643 7899 10646
rect 11973 10706 12039 10709
rect 12198 10706 12204 10708
rect 11973 10704 12204 10706
rect 11973 10648 11978 10704
rect 12034 10648 12204 10704
rect 11973 10646 12204 10648
rect 11973 10643 12039 10646
rect 12198 10644 12204 10646
rect 12268 10644 12274 10708
rect 5625 10570 5691 10573
rect 8109 10570 8175 10573
rect 10685 10570 10751 10573
rect 5625 10568 10751 10570
rect 5625 10512 5630 10568
rect 5686 10512 8114 10568
rect 8170 10512 10690 10568
rect 10746 10512 10751 10568
rect 5625 10510 10751 10512
rect 5625 10507 5691 10510
rect 8109 10507 8175 10510
rect 10685 10507 10751 10510
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 3785 10162 3851 10165
rect 8293 10162 8359 10165
rect 11329 10162 11395 10165
rect 3785 10160 11395 10162
rect 3785 10104 3790 10160
rect 3846 10104 8298 10160
rect 8354 10104 11334 10160
rect 11390 10104 11395 10160
rect 3785 10102 11395 10104
rect 3785 10099 3851 10102
rect 8293 10099 8359 10102
rect 11329 10099 11395 10102
rect 5257 10026 5323 10029
rect 9949 10026 10015 10029
rect 5257 10024 10015 10026
rect 5257 9968 5262 10024
rect 5318 9968 9954 10024
rect 10010 9968 10015 10024
rect 5257 9966 10015 9968
rect 5257 9963 5323 9966
rect 9949 9963 10015 9966
rect 8385 9890 8451 9893
rect 9305 9890 9371 9893
rect 8385 9888 9371 9890
rect 8385 9832 8390 9888
rect 8446 9832 9310 9888
rect 9366 9832 9371 9888
rect 8385 9830 9371 9832
rect 8385 9827 8451 9830
rect 9305 9827 9371 9830
rect 4906 9824 5302 9825
rect 4906 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5302 9824
rect 4906 9759 5302 9760
rect 10906 9824 11302 9825
rect 10906 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11302 9824
rect 10906 9759 11302 9760
rect 7189 9754 7255 9757
rect 8201 9754 8267 9757
rect 7189 9752 8267 9754
rect 7189 9696 7194 9752
rect 7250 9696 8206 9752
rect 8262 9696 8267 9752
rect 7189 9694 8267 9696
rect 7189 9691 7255 9694
rect 8201 9691 8267 9694
rect 3601 9618 3667 9621
rect 4889 9618 4955 9621
rect 3601 9616 4955 9618
rect 3601 9560 3606 9616
rect 3662 9560 4894 9616
rect 4950 9560 4955 9616
rect 3601 9558 4955 9560
rect 3601 9555 3667 9558
rect 4889 9555 4955 9558
rect 7005 9618 7071 9621
rect 8661 9618 8727 9621
rect 10777 9620 10843 9621
rect 10726 9618 10732 9620
rect 7005 9616 8727 9618
rect 7005 9560 7010 9616
rect 7066 9560 8666 9616
rect 8722 9560 8727 9616
rect 7005 9558 8727 9560
rect 10686 9558 10732 9618
rect 10796 9618 10843 9620
rect 10961 9618 11027 9621
rect 10796 9616 11027 9618
rect 10838 9560 10966 9616
rect 11022 9560 11027 9616
rect 7005 9555 7071 9558
rect 8661 9555 8727 9558
rect 10726 9556 10732 9558
rect 10796 9558 11027 9560
rect 10796 9556 10843 9558
rect 10777 9555 10843 9556
rect 10961 9555 11027 9558
rect 4613 9482 4679 9485
rect 6821 9482 6887 9485
rect 4613 9480 6887 9482
rect 4613 9424 4618 9480
rect 4674 9424 6826 9480
rect 6882 9424 6887 9480
rect 4613 9422 6887 9424
rect 4613 9419 4679 9422
rect 6821 9419 6887 9422
rect 8109 9482 8175 9485
rect 8753 9482 8819 9485
rect 8109 9480 8819 9482
rect 8109 9424 8114 9480
rect 8170 9424 8758 9480
rect 8814 9424 8819 9480
rect 8109 9422 8819 9424
rect 8109 9419 8175 9422
rect 8753 9419 8819 9422
rect 10685 9482 10751 9485
rect 10961 9482 11027 9485
rect 10685 9480 11027 9482
rect 10685 9424 10690 9480
rect 10746 9424 10966 9480
rect 11022 9424 11027 9480
rect 10685 9422 11027 9424
rect 10685 9419 10751 9422
rect 10961 9419 11027 9422
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 2313 9074 2379 9077
rect 5073 9074 5139 9077
rect 2313 9072 5139 9074
rect 2313 9016 2318 9072
rect 2374 9016 5078 9072
rect 5134 9016 5139 9072
rect 2313 9014 5139 9016
rect 2313 9011 2379 9014
rect 5073 9011 5139 9014
rect 6729 9074 6795 9077
rect 8569 9074 8635 9077
rect 6729 9072 8635 9074
rect 6729 9016 6734 9072
rect 6790 9016 8574 9072
rect 8630 9016 8635 9072
rect 6729 9014 8635 9016
rect 6729 9011 6795 9014
rect 8569 9011 8635 9014
rect 4981 8938 5047 8941
rect 7097 8938 7163 8941
rect 4981 8936 7163 8938
rect 4981 8880 4986 8936
rect 5042 8880 7102 8936
rect 7158 8880 7163 8936
rect 4981 8878 7163 8880
rect 4981 8875 5047 8878
rect 7097 8875 7163 8878
rect 4906 8736 5302 8737
rect 4906 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5302 8736
rect 4906 8671 5302 8672
rect 10906 8736 11302 8737
rect 10906 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11302 8736
rect 10906 8671 11302 8672
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 4906 7648 5302 7649
rect 4906 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5302 7648
rect 4906 7583 5302 7584
rect 10906 7648 11302 7649
rect 10906 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11302 7648
rect 10906 7583 11302 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 8477 7034 8543 7037
rect 9397 7034 9463 7037
rect 8477 7032 9463 7034
rect 8477 6976 8482 7032
rect 8538 6976 9402 7032
rect 9458 6976 9463 7032
rect 8477 6974 9463 6976
rect 8477 6971 8543 6974
rect 9397 6971 9463 6974
rect 8201 6762 8267 6765
rect 10685 6762 10751 6765
rect 8201 6760 10751 6762
rect 8201 6704 8206 6760
rect 8262 6704 10690 6760
rect 10746 6704 10751 6760
rect 8201 6702 10751 6704
rect 8201 6699 8267 6702
rect 10685 6699 10751 6702
rect 4906 6560 5302 6561
rect 4906 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5302 6560
rect 4906 6495 5302 6496
rect 10906 6560 11302 6561
rect 10906 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11302 6560
rect 10906 6495 11302 6496
rect 7005 6218 7071 6221
rect 7741 6218 7807 6221
rect 7005 6216 7807 6218
rect 7005 6160 7010 6216
rect 7066 6160 7746 6216
rect 7802 6160 7807 6216
rect 7005 6158 7807 6160
rect 7005 6155 7071 6158
rect 7741 6155 7807 6158
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 3233 5538 3299 5541
rect 3366 5538 3372 5540
rect 3233 5536 3372 5538
rect 3233 5480 3238 5536
rect 3294 5480 3372 5536
rect 3233 5478 3372 5480
rect 3233 5475 3299 5478
rect 3366 5476 3372 5478
rect 3436 5476 3442 5540
rect 4906 5472 5302 5473
rect 4906 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5302 5472
rect 4906 5407 5302 5408
rect 10906 5472 11302 5473
rect 10906 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11302 5472
rect 10906 5407 11302 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 4906 4384 5302 4385
rect 4906 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5302 4384
rect 4906 4319 5302 4320
rect 10906 4384 11302 4385
rect 10906 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11302 4384
rect 10906 4319 11302 4320
rect 3049 4042 3115 4045
rect 10317 4044 10383 4045
rect 3182 4042 3188 4044
rect 3049 4040 3188 4042
rect 3049 3984 3054 4040
rect 3110 3984 3188 4040
rect 3049 3982 3188 3984
rect 3049 3979 3115 3982
rect 3182 3980 3188 3982
rect 3252 3980 3258 4044
rect 10317 4042 10364 4044
rect 10272 4040 10364 4042
rect 10272 3984 10322 4040
rect 10272 3982 10364 3984
rect 10317 3980 10364 3982
rect 10428 3980 10434 4044
rect 10317 3979 10383 3980
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 4906 3296 5302 3297
rect 4906 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5302 3296
rect 4906 3231 5302 3232
rect 10906 3296 11302 3297
rect 10906 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11302 3296
rect 10906 3231 11302 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 4906 2208 5302 2209
rect 4906 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5302 2208
rect 4906 2143 5302 2144
rect 10906 2208 11302 2209
rect 10906 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11302 2208
rect 10906 2143 11302 2144
<< via3 >>
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 4912 14172 4976 14176
rect 4912 14116 4916 14172
rect 4916 14116 4972 14172
rect 4972 14116 4976 14172
rect 4912 14112 4976 14116
rect 4992 14172 5056 14176
rect 4992 14116 4996 14172
rect 4996 14116 5052 14172
rect 5052 14116 5056 14172
rect 4992 14112 5056 14116
rect 5072 14172 5136 14176
rect 5072 14116 5076 14172
rect 5076 14116 5132 14172
rect 5132 14116 5136 14172
rect 5072 14112 5136 14116
rect 5152 14172 5216 14176
rect 5152 14116 5156 14172
rect 5156 14116 5212 14172
rect 5212 14116 5216 14172
rect 5152 14112 5216 14116
rect 5232 14172 5296 14176
rect 5232 14116 5236 14172
rect 5236 14116 5292 14172
rect 5292 14116 5296 14172
rect 5232 14112 5296 14116
rect 10912 14172 10976 14176
rect 10912 14116 10916 14172
rect 10916 14116 10972 14172
rect 10972 14116 10976 14172
rect 10912 14112 10976 14116
rect 10992 14172 11056 14176
rect 10992 14116 10996 14172
rect 10996 14116 11052 14172
rect 11052 14116 11056 14172
rect 10992 14112 11056 14116
rect 11072 14172 11136 14176
rect 11072 14116 11076 14172
rect 11076 14116 11132 14172
rect 11132 14116 11136 14172
rect 11072 14112 11136 14116
rect 11152 14172 11216 14176
rect 11152 14116 11156 14172
rect 11156 14116 11212 14172
rect 11212 14116 11216 14172
rect 11152 14112 11216 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 10732 13772 10796 13836
rect 12204 13832 12268 13836
rect 12204 13776 12254 13832
rect 12254 13776 12268 13832
rect 12204 13772 12268 13776
rect 10364 13636 10428 13700
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 4912 13084 4976 13088
rect 4912 13028 4916 13084
rect 4916 13028 4972 13084
rect 4972 13028 4976 13084
rect 4912 13024 4976 13028
rect 4992 13084 5056 13088
rect 4992 13028 4996 13084
rect 4996 13028 5052 13084
rect 5052 13028 5056 13084
rect 4992 13024 5056 13028
rect 5072 13084 5136 13088
rect 5072 13028 5076 13084
rect 5076 13028 5132 13084
rect 5132 13028 5136 13084
rect 5072 13024 5136 13028
rect 5152 13084 5216 13088
rect 5152 13028 5156 13084
rect 5156 13028 5212 13084
rect 5212 13028 5216 13084
rect 5152 13024 5216 13028
rect 5232 13084 5296 13088
rect 5232 13028 5236 13084
rect 5236 13028 5292 13084
rect 5292 13028 5296 13084
rect 5232 13024 5296 13028
rect 10912 13084 10976 13088
rect 10912 13028 10916 13084
rect 10916 13028 10972 13084
rect 10972 13028 10976 13084
rect 10912 13024 10976 13028
rect 10992 13084 11056 13088
rect 10992 13028 10996 13084
rect 10996 13028 11052 13084
rect 11052 13028 11056 13084
rect 10992 13024 11056 13028
rect 11072 13084 11136 13088
rect 11072 13028 11076 13084
rect 11076 13028 11132 13084
rect 11132 13028 11136 13084
rect 11072 13024 11136 13028
rect 11152 13084 11216 13088
rect 11152 13028 11156 13084
rect 11156 13028 11212 13084
rect 11212 13028 11216 13084
rect 11152 13024 11216 13028
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 4912 11996 4976 12000
rect 4912 11940 4916 11996
rect 4916 11940 4972 11996
rect 4972 11940 4976 11996
rect 4912 11936 4976 11940
rect 4992 11996 5056 12000
rect 4992 11940 4996 11996
rect 4996 11940 5052 11996
rect 5052 11940 5056 11996
rect 4992 11936 5056 11940
rect 5072 11996 5136 12000
rect 5072 11940 5076 11996
rect 5076 11940 5132 11996
rect 5132 11940 5136 11996
rect 5072 11936 5136 11940
rect 5152 11996 5216 12000
rect 5152 11940 5156 11996
rect 5156 11940 5212 11996
rect 5212 11940 5216 11996
rect 5152 11936 5216 11940
rect 5232 11996 5296 12000
rect 5232 11940 5236 11996
rect 5236 11940 5292 11996
rect 5292 11940 5296 11996
rect 5232 11936 5296 11940
rect 10912 11996 10976 12000
rect 10912 11940 10916 11996
rect 10916 11940 10972 11996
rect 10972 11940 10976 11996
rect 10912 11936 10976 11940
rect 10992 11996 11056 12000
rect 10992 11940 10996 11996
rect 10996 11940 11052 11996
rect 11052 11940 11056 11996
rect 10992 11936 11056 11940
rect 11072 11996 11136 12000
rect 11072 11940 11076 11996
rect 11076 11940 11132 11996
rect 11132 11940 11136 11996
rect 11072 11936 11136 11940
rect 11152 11996 11216 12000
rect 11152 11940 11156 11996
rect 11156 11940 11212 11996
rect 11212 11940 11216 11996
rect 11152 11936 11216 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 3372 11248 3436 11252
rect 3372 11192 3422 11248
rect 3422 11192 3436 11248
rect 3372 11188 3436 11192
rect 3188 11112 3252 11116
rect 3188 11056 3238 11112
rect 3238 11056 3252 11112
rect 3188 11052 3252 11056
rect 4912 10908 4976 10912
rect 4912 10852 4916 10908
rect 4916 10852 4972 10908
rect 4972 10852 4976 10908
rect 4912 10848 4976 10852
rect 4992 10908 5056 10912
rect 4992 10852 4996 10908
rect 4996 10852 5052 10908
rect 5052 10852 5056 10908
rect 4992 10848 5056 10852
rect 5072 10908 5136 10912
rect 5072 10852 5076 10908
rect 5076 10852 5132 10908
rect 5132 10852 5136 10908
rect 5072 10848 5136 10852
rect 5152 10908 5216 10912
rect 5152 10852 5156 10908
rect 5156 10852 5212 10908
rect 5212 10852 5216 10908
rect 5152 10848 5216 10852
rect 5232 10908 5296 10912
rect 5232 10852 5236 10908
rect 5236 10852 5292 10908
rect 5292 10852 5296 10908
rect 5232 10848 5296 10852
rect 10912 10908 10976 10912
rect 10912 10852 10916 10908
rect 10916 10852 10972 10908
rect 10972 10852 10976 10908
rect 10912 10848 10976 10852
rect 10992 10908 11056 10912
rect 10992 10852 10996 10908
rect 10996 10852 11052 10908
rect 11052 10852 11056 10908
rect 10992 10848 11056 10852
rect 11072 10908 11136 10912
rect 11072 10852 11076 10908
rect 11076 10852 11132 10908
rect 11132 10852 11136 10908
rect 11072 10848 11136 10852
rect 11152 10908 11216 10912
rect 11152 10852 11156 10908
rect 11156 10852 11212 10908
rect 11212 10852 11216 10908
rect 11152 10848 11216 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 12204 10644 12268 10708
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 4912 9820 4976 9824
rect 4912 9764 4916 9820
rect 4916 9764 4972 9820
rect 4972 9764 4976 9820
rect 4912 9760 4976 9764
rect 4992 9820 5056 9824
rect 4992 9764 4996 9820
rect 4996 9764 5052 9820
rect 5052 9764 5056 9820
rect 4992 9760 5056 9764
rect 5072 9820 5136 9824
rect 5072 9764 5076 9820
rect 5076 9764 5132 9820
rect 5132 9764 5136 9820
rect 5072 9760 5136 9764
rect 5152 9820 5216 9824
rect 5152 9764 5156 9820
rect 5156 9764 5212 9820
rect 5212 9764 5216 9820
rect 5152 9760 5216 9764
rect 5232 9820 5296 9824
rect 5232 9764 5236 9820
rect 5236 9764 5292 9820
rect 5292 9764 5296 9820
rect 5232 9760 5296 9764
rect 10912 9820 10976 9824
rect 10912 9764 10916 9820
rect 10916 9764 10972 9820
rect 10972 9764 10976 9820
rect 10912 9760 10976 9764
rect 10992 9820 11056 9824
rect 10992 9764 10996 9820
rect 10996 9764 11052 9820
rect 11052 9764 11056 9820
rect 10992 9760 11056 9764
rect 11072 9820 11136 9824
rect 11072 9764 11076 9820
rect 11076 9764 11132 9820
rect 11132 9764 11136 9820
rect 11072 9760 11136 9764
rect 11152 9820 11216 9824
rect 11152 9764 11156 9820
rect 11156 9764 11212 9820
rect 11212 9764 11216 9820
rect 11152 9760 11216 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 10732 9616 10796 9620
rect 10732 9560 10782 9616
rect 10782 9560 10796 9616
rect 10732 9556 10796 9560
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 4912 8732 4976 8736
rect 4912 8676 4916 8732
rect 4916 8676 4972 8732
rect 4972 8676 4976 8732
rect 4912 8672 4976 8676
rect 4992 8732 5056 8736
rect 4992 8676 4996 8732
rect 4996 8676 5052 8732
rect 5052 8676 5056 8732
rect 4992 8672 5056 8676
rect 5072 8732 5136 8736
rect 5072 8676 5076 8732
rect 5076 8676 5132 8732
rect 5132 8676 5136 8732
rect 5072 8672 5136 8676
rect 5152 8732 5216 8736
rect 5152 8676 5156 8732
rect 5156 8676 5212 8732
rect 5212 8676 5216 8732
rect 5152 8672 5216 8676
rect 5232 8732 5296 8736
rect 5232 8676 5236 8732
rect 5236 8676 5292 8732
rect 5292 8676 5296 8732
rect 5232 8672 5296 8676
rect 10912 8732 10976 8736
rect 10912 8676 10916 8732
rect 10916 8676 10972 8732
rect 10972 8676 10976 8732
rect 10912 8672 10976 8676
rect 10992 8732 11056 8736
rect 10992 8676 10996 8732
rect 10996 8676 11052 8732
rect 11052 8676 11056 8732
rect 10992 8672 11056 8676
rect 11072 8732 11136 8736
rect 11072 8676 11076 8732
rect 11076 8676 11132 8732
rect 11132 8676 11136 8732
rect 11072 8672 11136 8676
rect 11152 8732 11216 8736
rect 11152 8676 11156 8732
rect 11156 8676 11212 8732
rect 11212 8676 11216 8732
rect 11152 8672 11216 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 4912 7644 4976 7648
rect 4912 7588 4916 7644
rect 4916 7588 4972 7644
rect 4972 7588 4976 7644
rect 4912 7584 4976 7588
rect 4992 7644 5056 7648
rect 4992 7588 4996 7644
rect 4996 7588 5052 7644
rect 5052 7588 5056 7644
rect 4992 7584 5056 7588
rect 5072 7644 5136 7648
rect 5072 7588 5076 7644
rect 5076 7588 5132 7644
rect 5132 7588 5136 7644
rect 5072 7584 5136 7588
rect 5152 7644 5216 7648
rect 5152 7588 5156 7644
rect 5156 7588 5212 7644
rect 5212 7588 5216 7644
rect 5152 7584 5216 7588
rect 5232 7644 5296 7648
rect 5232 7588 5236 7644
rect 5236 7588 5292 7644
rect 5292 7588 5296 7644
rect 5232 7584 5296 7588
rect 10912 7644 10976 7648
rect 10912 7588 10916 7644
rect 10916 7588 10972 7644
rect 10972 7588 10976 7644
rect 10912 7584 10976 7588
rect 10992 7644 11056 7648
rect 10992 7588 10996 7644
rect 10996 7588 11052 7644
rect 11052 7588 11056 7644
rect 10992 7584 11056 7588
rect 11072 7644 11136 7648
rect 11072 7588 11076 7644
rect 11076 7588 11132 7644
rect 11132 7588 11136 7644
rect 11072 7584 11136 7588
rect 11152 7644 11216 7648
rect 11152 7588 11156 7644
rect 11156 7588 11212 7644
rect 11212 7588 11216 7644
rect 11152 7584 11216 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 4912 6556 4976 6560
rect 4912 6500 4916 6556
rect 4916 6500 4972 6556
rect 4972 6500 4976 6556
rect 4912 6496 4976 6500
rect 4992 6556 5056 6560
rect 4992 6500 4996 6556
rect 4996 6500 5052 6556
rect 5052 6500 5056 6556
rect 4992 6496 5056 6500
rect 5072 6556 5136 6560
rect 5072 6500 5076 6556
rect 5076 6500 5132 6556
rect 5132 6500 5136 6556
rect 5072 6496 5136 6500
rect 5152 6556 5216 6560
rect 5152 6500 5156 6556
rect 5156 6500 5212 6556
rect 5212 6500 5216 6556
rect 5152 6496 5216 6500
rect 5232 6556 5296 6560
rect 5232 6500 5236 6556
rect 5236 6500 5292 6556
rect 5292 6500 5296 6556
rect 5232 6496 5296 6500
rect 10912 6556 10976 6560
rect 10912 6500 10916 6556
rect 10916 6500 10972 6556
rect 10972 6500 10976 6556
rect 10912 6496 10976 6500
rect 10992 6556 11056 6560
rect 10992 6500 10996 6556
rect 10996 6500 11052 6556
rect 11052 6500 11056 6556
rect 10992 6496 11056 6500
rect 11072 6556 11136 6560
rect 11072 6500 11076 6556
rect 11076 6500 11132 6556
rect 11132 6500 11136 6556
rect 11072 6496 11136 6500
rect 11152 6556 11216 6560
rect 11152 6500 11156 6556
rect 11156 6500 11212 6556
rect 11212 6500 11216 6556
rect 11152 6496 11216 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 3372 5476 3436 5540
rect 4912 5468 4976 5472
rect 4912 5412 4916 5468
rect 4916 5412 4972 5468
rect 4972 5412 4976 5468
rect 4912 5408 4976 5412
rect 4992 5468 5056 5472
rect 4992 5412 4996 5468
rect 4996 5412 5052 5468
rect 5052 5412 5056 5468
rect 4992 5408 5056 5412
rect 5072 5468 5136 5472
rect 5072 5412 5076 5468
rect 5076 5412 5132 5468
rect 5132 5412 5136 5468
rect 5072 5408 5136 5412
rect 5152 5468 5216 5472
rect 5152 5412 5156 5468
rect 5156 5412 5212 5468
rect 5212 5412 5216 5468
rect 5152 5408 5216 5412
rect 5232 5468 5296 5472
rect 5232 5412 5236 5468
rect 5236 5412 5292 5468
rect 5292 5412 5296 5468
rect 5232 5408 5296 5412
rect 10912 5468 10976 5472
rect 10912 5412 10916 5468
rect 10916 5412 10972 5468
rect 10972 5412 10976 5468
rect 10912 5408 10976 5412
rect 10992 5468 11056 5472
rect 10992 5412 10996 5468
rect 10996 5412 11052 5468
rect 11052 5412 11056 5468
rect 10992 5408 11056 5412
rect 11072 5468 11136 5472
rect 11072 5412 11076 5468
rect 11076 5412 11132 5468
rect 11132 5412 11136 5468
rect 11072 5408 11136 5412
rect 11152 5468 11216 5472
rect 11152 5412 11156 5468
rect 11156 5412 11212 5468
rect 11212 5412 11216 5468
rect 11152 5408 11216 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 4912 4380 4976 4384
rect 4912 4324 4916 4380
rect 4916 4324 4972 4380
rect 4972 4324 4976 4380
rect 4912 4320 4976 4324
rect 4992 4380 5056 4384
rect 4992 4324 4996 4380
rect 4996 4324 5052 4380
rect 5052 4324 5056 4380
rect 4992 4320 5056 4324
rect 5072 4380 5136 4384
rect 5072 4324 5076 4380
rect 5076 4324 5132 4380
rect 5132 4324 5136 4380
rect 5072 4320 5136 4324
rect 5152 4380 5216 4384
rect 5152 4324 5156 4380
rect 5156 4324 5212 4380
rect 5212 4324 5216 4380
rect 5152 4320 5216 4324
rect 5232 4380 5296 4384
rect 5232 4324 5236 4380
rect 5236 4324 5292 4380
rect 5292 4324 5296 4380
rect 5232 4320 5296 4324
rect 10912 4380 10976 4384
rect 10912 4324 10916 4380
rect 10916 4324 10972 4380
rect 10972 4324 10976 4380
rect 10912 4320 10976 4324
rect 10992 4380 11056 4384
rect 10992 4324 10996 4380
rect 10996 4324 11052 4380
rect 11052 4324 11056 4380
rect 10992 4320 11056 4324
rect 11072 4380 11136 4384
rect 11072 4324 11076 4380
rect 11076 4324 11132 4380
rect 11132 4324 11136 4380
rect 11072 4320 11136 4324
rect 11152 4380 11216 4384
rect 11152 4324 11156 4380
rect 11156 4324 11212 4380
rect 11212 4324 11216 4380
rect 11152 4320 11216 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 3188 3980 3252 4044
rect 10364 4040 10428 4044
rect 10364 3984 10378 4040
rect 10378 3984 10428 4040
rect 10364 3980 10428 3984
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 4912 3292 4976 3296
rect 4912 3236 4916 3292
rect 4916 3236 4972 3292
rect 4972 3236 4976 3292
rect 4912 3232 4976 3236
rect 4992 3292 5056 3296
rect 4992 3236 4996 3292
rect 4996 3236 5052 3292
rect 5052 3236 5056 3292
rect 4992 3232 5056 3236
rect 5072 3292 5136 3296
rect 5072 3236 5076 3292
rect 5076 3236 5132 3292
rect 5132 3236 5136 3292
rect 5072 3232 5136 3236
rect 5152 3292 5216 3296
rect 5152 3236 5156 3292
rect 5156 3236 5212 3292
rect 5212 3236 5216 3292
rect 5152 3232 5216 3236
rect 5232 3292 5296 3296
rect 5232 3236 5236 3292
rect 5236 3236 5292 3292
rect 5292 3236 5296 3292
rect 5232 3232 5296 3236
rect 10912 3292 10976 3296
rect 10912 3236 10916 3292
rect 10916 3236 10972 3292
rect 10972 3236 10976 3292
rect 10912 3232 10976 3236
rect 10992 3292 11056 3296
rect 10992 3236 10996 3292
rect 10996 3236 11052 3292
rect 11052 3236 11056 3292
rect 10992 3232 11056 3236
rect 11072 3292 11136 3296
rect 11072 3236 11076 3292
rect 11076 3236 11132 3292
rect 11132 3236 11136 3292
rect 11072 3232 11136 3236
rect 11152 3292 11216 3296
rect 11152 3236 11156 3292
rect 11156 3236 11212 3292
rect 11212 3236 11216 3292
rect 11152 3232 11216 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 4912 2204 4976 2208
rect 4912 2148 4916 2204
rect 4916 2148 4972 2204
rect 4972 2148 4976 2204
rect 4912 2144 4976 2148
rect 4992 2204 5056 2208
rect 4992 2148 4996 2204
rect 4996 2148 5052 2204
rect 5052 2148 5056 2204
rect 4992 2144 5056 2148
rect 5072 2204 5136 2208
rect 5072 2148 5076 2204
rect 5076 2148 5132 2204
rect 5132 2148 5136 2204
rect 5072 2144 5136 2148
rect 5152 2204 5216 2208
rect 5152 2148 5156 2204
rect 5156 2148 5212 2204
rect 5212 2148 5216 2204
rect 5152 2144 5216 2148
rect 5232 2204 5296 2208
rect 5232 2148 5236 2204
rect 5236 2148 5292 2204
rect 5292 2148 5296 2204
rect 5232 2144 5296 2148
rect 10912 2204 10976 2208
rect 10912 2148 10916 2204
rect 10916 2148 10972 2204
rect 10972 2148 10976 2204
rect 10912 2144 10976 2148
rect 10992 2204 11056 2208
rect 10992 2148 10996 2204
rect 10996 2148 11052 2204
rect 11052 2148 11056 2204
rect 10992 2144 11056 2148
rect 11072 2204 11136 2208
rect 11072 2148 11076 2204
rect 11076 2148 11132 2204
rect 11132 2148 11136 2204
rect 11072 2144 11136 2148
rect 11152 2204 11216 2208
rect 11152 2148 11156 2204
rect 11156 2148 11212 2204
rect 11212 2148 11216 2204
rect 11152 2144 11216 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
<< metal4 >>
rect 1904 14720 2304 14736
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 4904 14176 5304 14736
rect 4904 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5072 14176
rect 5136 14112 5152 14176
rect 5216 14112 5232 14176
rect 5296 14112 5304 14176
rect 4904 13088 5304 14112
rect 4904 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5072 13088
rect 5136 13024 5152 13088
rect 5216 13024 5232 13088
rect 5296 13024 5304 13088
rect 4904 12000 5304 13024
rect 4904 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5072 12000
rect 5136 11936 5152 12000
rect 5216 11936 5232 12000
rect 5296 11936 5304 12000
rect 3371 11252 3437 11253
rect 3371 11188 3372 11252
rect 3436 11188 3437 11252
rect 3371 11187 3437 11188
rect 3187 11116 3253 11117
rect 3187 11052 3188 11116
rect 3252 11052 3253 11116
rect 3187 11051 3253 11052
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9280 2304 10304
rect 1904 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 8192 2304 9216
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 3190 4045 3250 11051
rect 3374 5541 3434 11187
rect 4904 10912 5304 11936
rect 4904 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5072 10912
rect 5136 10848 5152 10912
rect 5216 10848 5232 10912
rect 5296 10848 5304 10912
rect 4904 9824 5304 10848
rect 4904 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5072 9824
rect 5136 9760 5152 9824
rect 5216 9760 5232 9824
rect 5296 9760 5304 9824
rect 4904 8736 5304 9760
rect 4904 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5072 8736
rect 5136 8672 5152 8736
rect 5216 8672 5232 8736
rect 5296 8672 5304 8736
rect 4904 7648 5304 8672
rect 4904 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5072 7648
rect 5136 7584 5152 7648
rect 5216 7584 5232 7648
rect 5296 7584 5304 7648
rect 4904 6560 5304 7584
rect 4904 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5072 6560
rect 5136 6496 5152 6560
rect 5216 6496 5232 6560
rect 5296 6496 5304 6560
rect 3371 5540 3437 5541
rect 3371 5476 3372 5540
rect 3436 5476 3437 5540
rect 3371 5475 3437 5476
rect 4904 5472 5304 6496
rect 4904 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5072 5472
rect 5136 5408 5152 5472
rect 5216 5408 5232 5472
rect 5296 5408 5304 5472
rect 4904 4384 5304 5408
rect 4904 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5072 4384
rect 5136 4320 5152 4384
rect 5216 4320 5232 4384
rect 5296 4320 5304 4384
rect 3187 4044 3253 4045
rect 3187 3980 3188 4044
rect 3252 3980 3253 4044
rect 3187 3979 3253 3980
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 2752 2304 3776
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 4904 3296 5304 4320
rect 4904 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5072 3296
rect 5136 3232 5152 3296
rect 5216 3232 5232 3296
rect 5296 3232 5304 3296
rect 4904 2208 5304 3232
rect 4904 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5072 2208
rect 5136 2144 5152 2208
rect 5216 2144 5232 2208
rect 5296 2144 5304 2208
rect 4904 2128 5304 2144
rect 7904 14720 8304 14736
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 10904 14176 11304 14736
rect 10904 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11072 14176
rect 11136 14112 11152 14176
rect 11216 14112 11232 14176
rect 11296 14112 11304 14176
rect 10731 13836 10797 13837
rect 10731 13772 10732 13836
rect 10796 13772 10797 13836
rect 10731 13771 10797 13772
rect 10363 13700 10429 13701
rect 10363 13636 10364 13700
rect 10428 13636 10429 13700
rect 10363 13635 10429 13636
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9280 8304 10304
rect 7904 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 8192 8304 9216
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 10366 4045 10426 13635
rect 10734 9621 10794 13771
rect 10904 13088 11304 14112
rect 12203 13836 12269 13837
rect 12203 13772 12204 13836
rect 12268 13772 12269 13836
rect 12203 13771 12269 13772
rect 10904 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11072 13088
rect 11136 13024 11152 13088
rect 11216 13024 11232 13088
rect 11296 13024 11304 13088
rect 10904 12000 11304 13024
rect 10904 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11072 12000
rect 11136 11936 11152 12000
rect 11216 11936 11232 12000
rect 11296 11936 11304 12000
rect 10904 10912 11304 11936
rect 10904 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11072 10912
rect 11136 10848 11152 10912
rect 11216 10848 11232 10912
rect 11296 10848 11304 10912
rect 10904 9824 11304 10848
rect 12206 10709 12266 13771
rect 12203 10708 12269 10709
rect 12203 10644 12204 10708
rect 12268 10644 12269 10708
rect 12203 10643 12269 10644
rect 10904 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11072 9824
rect 11136 9760 11152 9824
rect 11216 9760 11232 9824
rect 11296 9760 11304 9824
rect 10731 9620 10797 9621
rect 10731 9556 10732 9620
rect 10796 9556 10797 9620
rect 10731 9555 10797 9556
rect 10904 8736 11304 9760
rect 10904 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11072 8736
rect 11136 8672 11152 8736
rect 11216 8672 11232 8736
rect 11296 8672 11304 8736
rect 10904 7648 11304 8672
rect 10904 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11072 7648
rect 11136 7584 11152 7648
rect 11216 7584 11232 7648
rect 11296 7584 11304 7648
rect 10904 6560 11304 7584
rect 10904 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11072 6560
rect 11136 6496 11152 6560
rect 11216 6496 11232 6560
rect 11296 6496 11304 6560
rect 10904 5472 11304 6496
rect 10904 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11072 5472
rect 11136 5408 11152 5472
rect 11216 5408 11232 5472
rect 11296 5408 11304 5472
rect 10904 4384 11304 5408
rect 10904 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11072 4384
rect 11136 4320 11152 4384
rect 11216 4320 11232 4384
rect 11296 4320 11304 4384
rect 10363 4044 10429 4045
rect 10363 3980 10364 4044
rect 10428 3980 10429 4044
rect 10363 3979 10429 3980
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 2752 8304 3776
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 10904 3296 11304 4320
rect 10904 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11072 3296
rect 11136 3232 11152 3296
rect 11216 3232 11232 3296
rect 11296 3232 11304 3296
rect 10904 2208 11304 3232
rect 10904 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11072 2208
rect 11136 2144 11152 2208
rect 11216 2144 11232 2208
rect 11296 2144 11304 2208
rect 10904 2128 11304 2144
use sky130_fd_sc_hd__buf_2  _177_
timestamp 1713490400
transform 1 0 13248 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _178_
timestamp 1713490400
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _179_
timestamp 1713490400
transform -1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _180_
timestamp 1713490400
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 1713490400
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _182_
timestamp 1713490400
transform -1 0 9384 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _183_
timestamp 1713490400
transform -1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1713490400
transform -1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1713490400
transform 1 0 10212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_4  _186_
timestamp 1713490400
transform 1 0 11500 0 -1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_1  _187_
timestamp 1713490400
transform 1 0 8924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _188_
timestamp 1713490400
transform -1 0 9476 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1713490400
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _190_
timestamp 1713490400
transform -1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1713490400
transform -1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _192_
timestamp 1713490400
transform -1 0 8004 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _193_
timestamp 1713490400
transform -1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _194_
timestamp 1713490400
transform -1 0 11408 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1713490400
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o32ai_1  _196_
timestamp 1713490400
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _197_
timestamp 1713490400
transform 1 0 7268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _198_
timestamp 1713490400
transform -1 0 11408 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _199_
timestamp 1713490400
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _200_
timestamp 1713490400
transform 1 0 10764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _201_
timestamp 1713490400
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _202_
timestamp 1713490400
transform -1 0 11960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _203_
timestamp 1713490400
transform -1 0 11408 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _204_
timestamp 1713490400
transform -1 0 12236 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _205_
timestamp 1713490400
transform -1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _206_
timestamp 1713490400
transform -1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _207_
timestamp 1713490400
transform -1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _208_
timestamp 1713490400
transform 1 0 10396 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _209_
timestamp 1713490400
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_2  _210_
timestamp 1713490400
transform 1 0 4508 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_2  _211_
timestamp 1713490400
transform -1 0 10212 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 1713490400
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _213_
timestamp 1713490400
transform -1 0 8464 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _214_
timestamp 1713490400
transform 1 0 6716 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _215_
timestamp 1713490400
transform -1 0 9844 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_2  _216_
timestamp 1713490400
transform 1 0 7636 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _217_
timestamp 1713490400
transform -1 0 4508 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _218_
timestamp 1713490400
transform 1 0 4232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _219_
timestamp 1713490400
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _220_
timestamp 1713490400
transform -1 0 7544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _221_
timestamp 1713490400
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _222_
timestamp 1713490400
transform -1 0 3312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1713490400
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _224_
timestamp 1713490400
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _225_
timestamp 1713490400
transform -1 0 8924 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _226_
timestamp 1713490400
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _227_
timestamp 1713490400
transform -1 0 8004 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _228_
timestamp 1713490400
transform 1 0 6900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _229_
timestamp 1713490400
transform 1 0 2760 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _230_
timestamp 1713490400
transform 1 0 2944 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _231_
timestamp 1713490400
transform -1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1713490400
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _233_
timestamp 1713490400
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _234_
timestamp 1713490400
transform -1 0 8648 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _235_
timestamp 1713490400
transform 1 0 5796 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_2  _236_
timestamp 1713490400
transform 1 0 6348 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp 1713490400
transform -1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp 1713490400
transform -1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _239_
timestamp 1713490400
transform -1 0 10948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _240_
timestamp 1713490400
transform -1 0 10304 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _241_
timestamp 1713490400
transform -1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _242_
timestamp 1713490400
transform 1 0 6348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _243_
timestamp 1713490400
transform 1 0 9016 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _244_
timestamp 1713490400
transform 1 0 9844 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _245_
timestamp 1713490400
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _246_
timestamp 1713490400
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _247_
timestamp 1713490400
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _248_
timestamp 1713490400
transform -1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1713490400
transform -1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1713490400
transform -1 0 6900 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _251_
timestamp 1713490400
transform 1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _252_
timestamp 1713490400
transform 1 0 3956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _253_
timestamp 1713490400
transform -1 0 5336 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _254_
timestamp 1713490400
transform -1 0 5888 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1713490400
transform 1 0 4048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _256_
timestamp 1713490400
transform 1 0 4508 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _257_
timestamp 1713490400
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _258_
timestamp 1713490400
transform 1 0 4508 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _259_
timestamp 1713490400
transform -1 0 3772 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1713490400
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1713490400
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _262_
timestamp 1713490400
transform 1 0 8004 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _263_
timestamp 1713490400
transform -1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _264_
timestamp 1713490400
transform -1 0 8924 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _265_
timestamp 1713490400
transform -1 0 9660 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _266_
timestamp 1713490400
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _267_
timestamp 1713490400
transform -1 0 8280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1713490400
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1713490400
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _270_
timestamp 1713490400
transform 1 0 8280 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _271_
timestamp 1713490400
transform 1 0 10120 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1713490400
transform -1 0 7544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _273_
timestamp 1713490400
transform -1 0 7728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _274_
timestamp 1713490400
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _275_
timestamp 1713490400
transform -1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _276_
timestamp 1713490400
transform 1 0 3496 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _277_
timestamp 1713490400
transform -1 0 3496 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _278_
timestamp 1713490400
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_2  _279_
timestamp 1713490400
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1713490400
transform -1 0 8280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp 1713490400
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _282_
timestamp 1713490400
transform 1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _283_
timestamp 1713490400
transform -1 0 7728 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _284_
timestamp 1713490400
transform 1 0 11684 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _285_
timestamp 1713490400
transform -1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _286_
timestamp 1713490400
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _287_
timestamp 1713490400
transform 1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1713490400
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _289_
timestamp 1713490400
transform 1 0 8096 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1713490400
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _291_
timestamp 1713490400
transform 1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 1713490400
transform 1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1713490400
transform 1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _294_
timestamp 1713490400
transform 1 0 9660 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _295_
timestamp 1713490400
transform 1 0 9476 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _296_
timestamp 1713490400
transform 1 0 12788 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _297_
timestamp 1713490400
transform -1 0 12328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1713490400
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _299_
timestamp 1713490400
transform -1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp 1713490400
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _301_
timestamp 1713490400
transform 1 0 12144 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _302_
timestamp 1713490400
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _303_
timestamp 1713490400
transform 1 0 12328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _304_
timestamp 1713490400
transform 1 0 10672 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _305_
timestamp 1713490400
transform 1 0 11408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _306_
timestamp 1713490400
transform -1 0 11408 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _307_
timestamp 1713490400
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _308_
timestamp 1713490400
transform -1 0 8372 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _309_
timestamp 1713490400
transform -1 0 7360 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _310_
timestamp 1713490400
transform -1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _311_
timestamp 1713490400
transform -1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _312_
timestamp 1713490400
transform -1 0 6992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _313_
timestamp 1713490400
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _314_
timestamp 1713490400
transform 1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _315_
timestamp 1713490400
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _316_
timestamp 1713490400
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _317_
timestamp 1713490400
transform 1 0 3036 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _318_
timestamp 1713490400
transform 1 0 2760 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 1713490400
transform -1 0 4416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _320_
timestamp 1713490400
transform 1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _321_
timestamp 1713490400
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _322_
timestamp 1713490400
transform -1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _323_
timestamp 1713490400
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _324_
timestamp 1713490400
transform 1 0 4784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _325_
timestamp 1713490400
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _326_
timestamp 1713490400
transform -1 0 6164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _327_
timestamp 1713490400
transform -1 0 7728 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _328_
timestamp 1713490400
transform -1 0 5428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp 1713490400
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _330_
timestamp 1713490400
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _331_
timestamp 1713490400
transform -1 0 9752 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _332_
timestamp 1713490400
transform 1 0 8372 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _333_
timestamp 1713490400
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _334_
timestamp 1713490400
transform -1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _335_
timestamp 1713490400
transform 1 0 9476 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _336_
timestamp 1713490400
transform 1 0 10120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _337_
timestamp 1713490400
transform 1 0 6808 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _338_
timestamp 1713490400
transform -1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _339_
timestamp 1713490400
transform 1 0 11500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _340_
timestamp 1713490400
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _341_
timestamp 1713490400
transform 1 0 9844 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1713490400
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _343_
timestamp 1713490400
transform 1 0 10672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _344_
timestamp 1713490400
transform 1 0 10396 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _345_
timestamp 1713490400
transform 1 0 9752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _346_
timestamp 1713490400
transform -1 0 5336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _347_
timestamp 1713490400
transform 1 0 4600 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _348_
timestamp 1713490400
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _349_
timestamp 1713490400
transform -1 0 6256 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _350_
timestamp 1713490400
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _351_
timestamp 1713490400
transform 1 0 3864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _352_
timestamp 1713490400
transform 1 0 3312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1713490400
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 1713490400
transform 1 0 2024 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _355_
timestamp 1713490400
transform 1 0 1472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 1713490400
transform 1 0 2024 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _357_
timestamp 1713490400
transform 1 0 3956 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 1713490400
transform 1 0 2300 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _359_
timestamp 1713490400
transform -1 0 13616 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _360_
timestamp 1713490400
transform 1 0 7360 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _361_
timestamp 1713490400
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _362_
timestamp 1713490400
transform -1 0 6900 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 1713490400
transform -1 0 2944 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _364_
timestamp 1713490400
transform 1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1713490400
transform -1 0 10396 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _366_
timestamp 1713490400
transform -1 0 11868 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _367_
timestamp 1713490400
transform 1 0 12144 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1713490400
transform 1 0 11868 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1713490400
transform -1 0 2944 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1713490400
transform 1 0 1564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1713490400
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1713490400
transform 1 0 3496 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1713490400
transform 1 0 4600 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1713490400
transform 1 0 4416 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1713490400
transform 1 0 5888 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1713490400
transform 1 0 5428 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1713490400
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1713490400
transform 1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _379_
timestamp 1713490400
transform 1 0 6164 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1713490400
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1713490400
transform 1 0 10396 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1713490400
transform 1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1713490400
transform 1 0 4048 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1713490400
transform 1 0 2760 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1713490400
transform 1 0 12144 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1713490400
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1713490400
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1713490400
transform -1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1713490400
transform -1 0 6072 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1713490400
transform -1 0 6348 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1713490400
transform 1 0 10488 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1713490400
transform 1 0 10672 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6
timestamp 1713490400
transform 1 0 1656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_12
timestamp 1713490400
transform 1 0 2208 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16
timestamp 1713490400
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_32
timestamp 1713490400
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_38
timestamp 1713490400
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_48
timestamp 1713490400
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1713490400
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1713490400
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_68
timestamp 1713490400
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_76
timestamp 1713490400
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1713490400
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85
timestamp 1713490400
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_94
timestamp 1713490400
transform 1 0 9752 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_102
timestamp 1713490400
transform 1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_107
timestamp 1713490400
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1713490400
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1713490400
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_120
timestamp 1713490400
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_128
timestamp 1713490400
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_133
timestamp 1713490400
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1713490400
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_15
timestamp 1713490400
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 1713490400
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_35
timestamp 1713490400
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1713490400
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_63
timestamp 1713490400
transform 1 0 6900 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_75
timestamp 1713490400
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_79
timestamp 1713490400
transform 1 0 8372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_87
timestamp 1713490400
transform 1 0 9108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_97
timestamp 1713490400
transform 1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102
timestamp 1713490400
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1713490400
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1713490400
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1713490400
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_137
timestamp 1713490400
transform 1 0 13708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_3
timestamp 1713490400
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_11
timestamp 1713490400
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1713490400
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_117
timestamp 1713490400
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_129
timestamp 1713490400
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_137
timestamp 1713490400
transform 1 0 13708 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1713490400
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_15
timestamp 1713490400
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_42
timestamp 1713490400
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_46
timestamp 1713490400
transform 1 0 5336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1713490400
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_63
timestamp 1713490400
transform 1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_90
timestamp 1713490400
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_113
timestamp 1713490400
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1713490400
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_136
timestamp 1713490400
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1713490400
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1713490400
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1713490400
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp 1713490400
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_48
timestamp 1713490400
transform 1 0 5520 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_60
timestamp 1713490400
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_72
timestamp 1713490400
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1713490400
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_94
timestamp 1713490400
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_104
timestamp 1713490400
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_116
timestamp 1713490400
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_136
timestamp 1713490400
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1713490400
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_28
timestamp 1713490400
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1713490400
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1713490400
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1713490400
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 1713490400
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_73
timestamp 1713490400
transform 1 0 7820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_85
timestamp 1713490400
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_100
timestamp 1713490400
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1713490400
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_129
timestamp 1713490400
transform 1 0 12972 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_137
timestamp 1713490400
transform 1 0 13708 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_3
timestamp 1713490400
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1713490400
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_35
timestamp 1713490400
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_68
timestamp 1713490400
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_80
timestamp 1713490400
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_92
timestamp 1713490400
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_122
timestamp 1713490400
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_134
timestamp 1713490400
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1713490400
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_9
timestamp 1713490400
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1713490400
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1713490400
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_72
timestamp 1713490400
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_93
timestamp 1713490400
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1713490400
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1713490400
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_137
timestamp 1713490400
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1713490400
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1713490400
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1713490400
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 1713490400
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_48
timestamp 1713490400
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_72
timestamp 1713490400
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_90
timestamp 1713490400
transform 1 0 9384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_96
timestamp 1713490400
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_104
timestamp 1713490400
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_132
timestamp 1713490400
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1713490400
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1713490400
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 1713490400
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_41
timestamp 1713490400
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1713490400
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1713490400
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1713490400
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_68
timestamp 1713490400
transform 1 0 7360 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_76
timestamp 1713490400
transform 1 0 8096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_92
timestamp 1713490400
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 1713490400
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1713490400
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_15
timestamp 1713490400
transform 1 0 2484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1713490400
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1713490400
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1713490400
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_43
timestamp 1713490400
transform 1 0 5060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_55
timestamp 1713490400
transform 1 0 6164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_67
timestamp 1713490400
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1713490400
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_90
timestamp 1713490400
transform 1 0 9384 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_98
timestamp 1713490400
transform 1 0 10120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_129
timestamp 1713490400
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_137
timestamp 1713490400
transform 1 0 13708 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1713490400
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1713490400
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 1713490400
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1713490400
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1713490400
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_67
timestamp 1713490400
transform 1 0 7268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_90
timestamp 1713490400
transform 1 0 9384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_98
timestamp 1713490400
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 1713490400
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1713490400
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_121
timestamp 1713490400
transform 1 0 12236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_128
timestamp 1713490400
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_136
timestamp 1713490400
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1713490400
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1713490400
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_56
timestamp 1713490400
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_75
timestamp 1713490400
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1713490400
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_92
timestamp 1713490400
transform 1 0 9568 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_100
timestamp 1713490400
transform 1 0 10304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_112
timestamp 1713490400
transform 1 0 11408 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_136
timestamp 1713490400
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1713490400
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_7
timestamp 1713490400
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_17
timestamp 1713490400
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_26
timestamp 1713490400
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_47
timestamp 1713490400
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1713490400
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_88
timestamp 1713490400
transform 1 0 9200 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_94
timestamp 1713490400
transform 1 0 9752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1713490400
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_121
timestamp 1713490400
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_133
timestamp 1713490400
transform 1 0 13340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_137
timestamp 1713490400
transform 1 0 13708 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1713490400
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1713490400
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1713490400
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1713490400
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1713490400
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1713490400
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_102
timestamp 1713490400
transform 1 0 10488 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_124
timestamp 1713490400
transform 1 0 12512 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_136
timestamp 1713490400
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1713490400
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_15
timestamp 1713490400
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_34
timestamp 1713490400
transform 1 0 4232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_38
timestamp 1713490400
transform 1 0 4600 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_47
timestamp 1713490400
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1713490400
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_66
timestamp 1713490400
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_81
timestamp 1713490400
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_85
timestamp 1713490400
transform 1 0 8924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_89
timestamp 1713490400
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1713490400
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1713490400
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_129
timestamp 1713490400
transform 1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_137
timestamp 1713490400
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1713490400
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1713490400
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 1713490400
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_43
timestamp 1713490400
transform 1 0 5060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_55
timestamp 1713490400
transform 1 0 6164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_61
timestamp 1713490400
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_65
timestamp 1713490400
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_69
timestamp 1713490400
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1713490400
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1713490400
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_102
timestamp 1713490400
transform 1 0 10488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_132
timestamp 1713490400
transform 1 0 13248 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1713490400
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_15
timestamp 1713490400
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_29
timestamp 1713490400
transform 1 0 3772 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1713490400
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1713490400
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1713490400
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_77
timestamp 1713490400
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_89
timestamp 1713490400
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_100
timestamp 1713490400
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_137
timestamp 1713490400
transform 1 0 13708 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1713490400
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_44
timestamp 1713490400
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_55
timestamp 1713490400
transform 1 0 6164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_63
timestamp 1713490400
transform 1 0 6900 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_70
timestamp 1713490400
transform 1 0 7544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1713490400
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1713490400
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_129
timestamp 1713490400
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_137
timestamp 1713490400
transform 1 0 13708 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_3
timestamp 1713490400
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_9
timestamp 1713490400
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_29
timestamp 1713490400
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1713490400
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1713490400
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_122
timestamp 1713490400
transform 1 0 12328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_134
timestamp 1713490400
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1713490400
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1713490400
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1713490400
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_29
timestamp 1713490400
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_63
timestamp 1713490400
transform 1 0 6900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1713490400
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1713490400
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_91
timestamp 1713490400
transform 1 0 9476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_99
timestamp 1713490400
transform 1 0 10212 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_133
timestamp 1713490400
transform 1 0 13340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_137
timestamp 1713490400
transform 1 0 13708 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1713490400
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_15
timestamp 1713490400
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_19
timestamp 1713490400
transform 1 0 2852 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_29
timestamp 1713490400
transform 1 0 3772 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_35
timestamp 1713490400
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1713490400
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1713490400
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_68
timestamp 1713490400
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_80
timestamp 1713490400
transform 1 0 8464 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1713490400
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1713490400
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1713490400
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_137
timestamp 1713490400
transform 1 0 13708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_6
timestamp 1713490400
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_10
timestamp 1713490400
transform 1 0 2024 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_14
timestamp 1713490400
transform 1 0 2392 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1713490400
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_29
timestamp 1713490400
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_36
timestamp 1713490400
transform 1 0 4416 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_47
timestamp 1713490400
transform 1 0 5428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_55
timestamp 1713490400
transform 1 0 6164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_60
timestamp 1713490400
transform 1 0 6624 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_69
timestamp 1713490400
transform 1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1713490400
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 1713490400
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_91
timestamp 1713490400
transform 1 0 9476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_103
timestamp 1713490400
transform 1 0 10580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_111
timestamp 1713490400
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_116
timestamp 1713490400
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_120
timestamp 1713490400
transform 1 0 12144 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_124
timestamp 1713490400
transform 1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_136
timestamp 1713490400
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1713490400
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1713490400
transform -1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1713490400
transform -1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1713490400
transform -1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1713490400
transform -1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1713490400
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1713490400
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1713490400
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1713490400
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 1713490400
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1713490400
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1713490400
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1713490400
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 1713490400
transform -1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 1713490400
transform -1 0 9476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1713490400
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1713490400
transform 1 0 7176 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 1713490400
transform -1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1713490400
transform 1 0 5152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1713490400
transform 1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1713490400
transform 1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output22
timestamp 1713490400
transform -1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1713490400
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output24
timestamp 1713490400
transform -1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 1713490400
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1713490400
transform -1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 1713490400
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1713490400
transform -1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 1713490400
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1713490400
transform -1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 1713490400
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1713490400
transform -1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 1713490400
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1713490400
transform -1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 1713490400
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1713490400
transform -1 0 14076 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 1713490400
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1713490400
transform -1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 1713490400
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1713490400
transform -1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 1713490400
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1713490400
transform -1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 1713490400
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1713490400
transform -1 0 14076 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 1713490400
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1713490400
transform -1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 1713490400
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1713490400
transform -1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 1713490400
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1713490400
transform -1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 1713490400
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1713490400
transform -1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 1713490400
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1713490400
transform -1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 1713490400
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1713490400
transform -1 0 14076 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 1713490400
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1713490400
transform -1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 1713490400
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1713490400
transform -1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 1713490400
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1713490400
transform -1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 1713490400
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1713490400
transform -1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 1713490400
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1713490400
transform -1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 1713490400
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1713490400
transform -1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 1713490400
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1713490400
transform -1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46
timestamp 1713490400
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 1713490400
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 1713490400
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 1713490400
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp 1713490400
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp 1713490400
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp 1713490400
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 1713490400
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp 1713490400
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp 1713490400
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp 1713490400
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp 1713490400
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 1713490400
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 1713490400
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp 1713490400
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp 1713490400
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1713490400
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1713490400
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_64
timestamp 1713490400
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 1713490400
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_66
timestamp 1713490400
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_67
timestamp 1713490400
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_68
timestamp 1713490400
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_69
timestamp 1713490400
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_70
timestamp 1713490400
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_71
timestamp 1713490400
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_72
timestamp 1713490400
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_73
timestamp 1713490400
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_74
timestamp 1713490400
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_75
timestamp 1713490400
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_76
timestamp 1713490400
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_77
timestamp 1713490400
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_78
timestamp 1713490400
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_79
timestamp 1713490400
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp 1713490400
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_81
timestamp 1713490400
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_82
timestamp 1713490400
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_83
timestamp 1713490400
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_84
timestamp 1713490400
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_85
timestamp 1713490400
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_86
timestamp 1713490400
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_87
timestamp 1713490400
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_88
timestamp 1713490400
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_89
timestamp 1713490400
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp 1713490400
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp 1713490400
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_92
timestamp 1713490400
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_93
timestamp 1713490400
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_94
timestamp 1713490400
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_95
timestamp 1713490400
transform 1 0 11408 0 1 14144
box -38 -48 130 592
<< labels >>
rlabel metal1 s 7590 14144 7590 14144 4 VGND
rlabel metal1 s 7590 14688 7590 14688 4 VPWR
rlabel metal1 s 2479 7446 2479 7446 4 _000_
rlabel metal2 s 1789 8874 1789 8874 4 _001_
rlabel metal1 s 2300 12954 2300 12954 4 _002_
rlabel metal1 s 4273 13294 4273 13294 4 _003_
rlabel metal2 s 2990 13260 2990 13260 4 _004_
rlabel metal1 s 7723 3434 7723 3434 4 _005_
rlabel metal1 s 9138 3434 9138 3434 4 _006_
rlabel metal1 s 6490 13226 6490 13226 4 _007_
rlabel metal1 s 2821 11050 2821 11050 4 _008_
rlabel metal2 s 7682 13090 7682 13090 4 _009_
rlabel metal1 s 9480 12818 9480 12818 4 _010_
rlabel metal1 s 10304 12410 10304 12410 4 _011_
rlabel metal1 s 12461 11730 12461 11730 4 _012_
rlabel metal1 s 12190 12886 12190 12886 4 _013_
rlabel metal1 s 2821 5270 2821 5270 4 _014_
rlabel metal1 s 1881 5678 1881 5678 4 _015_
rlabel metal1 s 2571 3434 2571 3434 4 _016_
rlabel metal1 s 3905 4182 3905 4182 4 _017_
rlabel metal1 s 4814 3094 4814 3094 4 _018_
rlabel metal1 s 4779 3434 4779 3434 4 _019_
rlabel metal2 s 6205 3502 6205 3502 4 _020_
rlabel metal1 s 5550 5610 5550 5610 4 _021_
rlabel metal1 s 11668 5270 11668 5270 4 _022_
rlabel metal1 s 11863 6698 11863 6698 4 _023_
rlabel metal1 s 6240 6698 6240 6698 4 _024_
rlabel metal1 s 12006 8976 12006 8976 4 _025_
rlabel metal2 s 10713 3502 10713 3502 4 _026_
rlabel metal1 s 10018 4114 10018 4114 4 _027_
rlabel metal2 s 4365 6766 4365 6766 4 _028_
rlabel metal1 s 3307 6358 3307 6358 4 _029_
rlabel metal1 s 8786 9894 8786 9894 4 _030_
rlabel metal1 s 4186 9675 4186 9675 4 _031_
rlabel metal1 s 6854 10438 6854 10438 4 _032_
rlabel metal1 s 8878 9588 8878 9588 4 _033_
rlabel metal1 s 4554 9962 4554 9962 4 _034_
rlabel metal1 s 4646 9486 4646 9486 4 _035_
rlabel metal1 s 11730 8908 11730 8908 4 _036_
rlabel metal1 s 3128 8534 3128 8534 4 _037_
rlabel metal1 s 7268 8874 7268 8874 4 _038_
rlabel metal1 s 3128 8330 3128 8330 4 _039_
rlabel metal2 s 2806 8058 2806 8058 4 _040_
rlabel metal1 s 4370 10642 4370 10642 4 _041_
rlabel metal1 s 7038 9962 7038 9962 4 _042_
rlabel metal1 s 3358 9452 3358 9452 4 _043_
rlabel metal1 s 7498 9146 7498 9146 4 _044_
rlabel metal1 s 3358 9554 3358 9554 4 _045_
rlabel metal1 s 2714 9486 2714 9486 4 _046_
rlabel metal2 s 2898 9656 2898 9656 4 _047_
rlabel metal1 s 2116 9554 2116 9554 4 _048_
rlabel metal1 s 8004 7242 8004 7242 4 _049_
rlabel metal1 s 4692 12954 4692 12954 4 _050_
rlabel metal1 s 6578 10098 6578 10098 4 _051_
rlabel metal1 s 4048 10642 4048 10642 4 _052_
rlabel metal1 s 6987 10982 6987 10982 4 _053_
rlabel metal1 s 4922 10506 4922 10506 4 _054_
rlabel metal1 s 10304 12614 10304 12614 4 _055_
rlabel metal1 s 11270 12852 11270 12852 4 _056_
rlabel metal1 s 8648 10506 8648 10506 4 _057_
rlabel metal1 s 5198 10676 5198 10676 4 _058_
rlabel metal2 s 10074 11729 10074 11729 4 _059_
rlabel metal1 s 10166 10098 10166 10098 4 _060_
rlabel metal1 s 3818 11662 3818 11662 4 _061_
rlabel metal1 s 3036 11866 3036 11866 4 _062_
rlabel metal1 s 2898 12342 2898 12342 4 _063_
rlabel metal1 s 2438 12410 2438 12410 4 _064_
rlabel metal1 s 6532 12410 6532 12410 4 _065_
rlabel metal1 s 5152 12750 5152 12750 4 _066_
rlabel metal1 s 5842 12682 5842 12682 4 _067_
rlabel metal1 s 5382 12682 5382 12682 4 _068_
rlabel metal2 s 5382 13430 5382 13430 4 _069_
rlabel metal1 s 4508 12206 4508 12206 4 _070_
rlabel metal1 s 3772 12410 3772 12410 4 _071_
rlabel metal1 s 4002 13770 4002 13770 4 _072_
rlabel metal1 s 3174 13872 3174 13872 4 _073_
rlabel metal1 s 9062 4114 9062 4114 4 _074_
rlabel metal1 s 6946 6290 6946 6290 4 _075_
rlabel metal1 s 9154 4794 9154 4794 4 _076_
rlabel metal1 s 7912 7310 7912 7310 4 _077_
rlabel metal1 s 9292 4114 9292 4114 4 _078_
rlabel metal1 s 8740 4114 8740 4114 4 _079_
rlabel metal2 s 8510 3502 8510 3502 4 _080_
rlabel metal1 s 10396 5678 10396 5678 4 _081_
rlabel metal1 s 7498 12240 7498 12240 4 _082_
rlabel metal1 s 7084 12410 7084 12410 4 _083_
rlabel metal2 s 7038 13362 7038 13362 4 _084_
rlabel metal3 s 8142 10557 8142 10557 4 _085_
rlabel metal1 s 3496 10778 3496 10778 4 _086_
rlabel metal1 s 3450 10608 3450 10608 4 _087_
rlabel metal1 s 8924 12750 8924 12750 4 _088_
rlabel metal1 s 6854 12818 6854 12818 4 _089_
rlabel metal1 s 7038 12954 7038 12954 4 _090_
rlabel metal1 s 7222 12886 7222 12886 4 _091_
rlabel metal1 s 11914 11662 11914 11662 4 _092_
rlabel metal2 s 8326 13022 8326 13022 4 _093_
rlabel metal1 s 7774 11798 7774 11798 4 _094_
rlabel metal1 s 7360 11866 7360 11866 4 _095_
rlabel metal1 s 8142 12410 8142 12410 4 _096_
rlabel metal1 s 11132 12614 11132 12614 4 _097_
rlabel metal1 s 8510 11084 8510 11084 4 _098_
rlabel metal1 s 10902 11866 10902 11866 4 _099_
rlabel metal1 s 10212 11662 10212 11662 4 _100_
rlabel metal1 s 9890 11866 9890 11866 4 _101_
rlabel metal2 s 13202 11424 13202 11424 4 _102_
rlabel metal1 s 11776 11730 11776 11730 4 _103_
rlabel metal1 s 11638 10744 11638 10744 4 _104_
rlabel metal1 s 12236 11866 12236 11866 4 _105_
rlabel metal2 s 10626 6052 10626 6052 4 _106_
rlabel metal1 s 12512 10574 12512 10574 4 _107_
rlabel metal2 s 12650 11492 12650 11492 4 _108_
rlabel metal1 s 11224 10778 11224 10778 4 _109_
rlabel metal1 s 11178 11186 11178 11186 4 _110_
rlabel metal1 s 11592 11322 11592 11322 4 _111_
rlabel metal1 s 8188 6154 8188 6154 4 _112_
rlabel metal1 s 6808 5202 6808 5202 4 _113_
rlabel metal1 s 2438 6324 2438 6324 4 _114_
rlabel metal2 s 9798 6766 9798 6766 4 _115_
rlabel metal1 s 6900 6154 6900 6154 4 _116_
rlabel metal1 s 3450 5236 3450 5236 4 _117_
rlabel metal2 s 2530 6086 2530 6086 4 _118_
rlabel metal1 s 3174 3162 3174 3162 4 _119_
rlabel metal1 s 4416 3706 4416 3706 4 _120_
rlabel metal1 s 4830 2618 4830 2618 4 _121_
rlabel metal2 s 6394 4386 6394 4386 4 _122_
rlabel metal1 s 6026 3162 6026 3162 4 _123_
rlabel metal1 s 4922 5644 4922 5644 4 _124_
rlabel metal1 s 10396 6970 10396 6970 4 _125_
rlabel metal1 s 10580 5134 10580 5134 4 _126_
rlabel metal2 s 9706 4998 9706 4998 4 _127_
rlabel metal1 s 9614 5236 9614 5236 4 _128_
rlabel metal1 s 9890 5168 9890 5168 4 _129_
rlabel metal1 s 10166 6834 10166 6834 4 _130_
rlabel metal2 s 6118 6970 6118 6970 4 _131_
rlabel metal1 s 10258 4658 10258 4658 4 _132_
rlabel metal1 s 11086 5202 11086 5202 4 _133_
rlabel metal1 s 10626 5236 10626 5236 4 _134_
rlabel metal1 s 10350 5338 10350 5338 4 _135_
rlabel metal1 s 4830 7888 4830 7888 4 _136_
rlabel metal1 s 4600 7854 4600 7854 4 _137_
rlabel metal2 s 4554 8772 4554 8772 4 _138_
rlabel metal1 s 3634 8398 3634 8398 4 _139_
rlabel metal1 s 3542 8330 3542 8330 4 _140_
rlabel metal1 s 3772 7378 3772 7378 4 _141_
rlabel metal2 s 8970 7616 8970 7616 4 _142_
rlabel metal1 s 9154 7310 9154 7310 4 _143_
rlabel metal1 s 8694 7786 8694 7786 4 _144_
rlabel metal1 s 8004 6970 8004 6970 4 _145_
rlabel metal2 s 9338 7378 9338 7378 4 _146_
rlabel metal1 s 8464 9146 8464 9146 4 _147_
rlabel metal2 s 7038 7820 7038 7820 4 _148_
rlabel metal1 s 8832 10642 8832 10642 4 _149_
rlabel metal2 s 9890 10880 9890 10880 4 _150_
rlabel metal2 s 8188 9350 8188 9350 4 _151_
rlabel metal1 s 7958 10132 7958 10132 4 _152_
rlabel metal1 s 5750 8976 5750 8976 4 _153_
rlabel metal2 s 7222 10574 7222 10574 4 _154_
rlabel metal1 s 7636 12818 7636 12818 4 _155_
rlabel metal2 s 7406 11628 7406 11628 4 _156_
rlabel metal1 s 4692 9554 4692 9554 4 _157_
rlabel metal1 s 11638 6426 11638 6426 4 _158_
rlabel metal1 s 9522 7412 9522 7412 4 _159_
rlabel metal1 s 10488 6222 10488 6222 4 _160_
rlabel metal1 s 7498 9996 7498 9996 4 _161_
rlabel metal1 s 6164 9690 6164 9690 4 _162_
rlabel metal1 s 10120 9554 10120 9554 4 _163_
rlabel metal1 s 9660 6290 9660 6290 4 _164_
rlabel metal1 s 10534 6902 10534 6902 4 _165_
rlabel metal2 s 10258 8534 10258 8534 4 _166_
rlabel metal1 s 8372 10030 8372 10030 4 _167_
rlabel metal1 s 10810 9078 10810 9078 4 _168_
rlabel metal2 s 10626 8432 10626 8432 4 _169_
rlabel metal1 s 12144 8058 12144 8058 4 _170_
rlabel metal1 s 12190 9520 12190 9520 4 _171_
rlabel metal1 s 8142 11628 8142 11628 4 _172_
rlabel metal2 s 10442 9350 10442 9350 4 _173_
rlabel metal3 s 7682 9044 7682 9044 4 _174_
rlabel metal1 s 4462 9690 4462 9690 4 _175_
rlabel metal2 s 9890 9452 9890 9452 4 _176_
rlabel metal1 s 13524 4250 13524 4250 4 adc.comparator.compres.ffsync.stage0
rlabel metal1 s 10442 4488 10442 4488 4 adc.comparator.compres.ffsync.stage1
rlabel metal1 s 9108 13498 9108 13498 4 adc.internalCounter\[0\]
rlabel metal1 s 10580 12886 10580 12886 4 adc.internalCounter\[1\]
rlabel metal1 s 9246 10608 9246 10608 4 adc.internalCounter\[2\]
rlabel metal1 s 12190 9622 12190 9622 4 adc.internalCounter\[3\]
rlabel metal1 s 9522 9996 9522 9996 4 adc.internalCounter\[4\]
rlabel metal1 s 12742 6290 12742 6290 4 adc.state\[0\]
rlabel metal2 s 12834 6426 12834 6426 4 adc.state\[1\]
rlabel metal1 s 8050 6732 8050 6732 4 adc.state\[2\]
rlabel metal1 s 13202 8466 13202 8466 4 adc.state\[3\]
rlabel metal1 s 8786 3094 8786 3094 4 adc.syncroCount\[0\]
rlabel metal2 s 8694 3298 8694 3298 4 adc.syncroCount\[1\]
rlabel metal2 s 14214 1588 14214 1588 4 analog_comparator_out
rlabel metal2 s 12190 15514 12190 15514 4 calib_enable
rlabel metal2 s 14214 12590 14214 12590 4 clk
rlabel metal1 s 10626 9962 10626 9962 4 clknet_0_clk
rlabel metal1 s 1610 5610 1610 5610 4 clknet_2_0__leaf_clk
rlabel metal1 s 2162 8942 2162 8942 4 clknet_2_1__leaf_clk
rlabel metal1 s 8188 3502 8188 3502 4 clknet_2_2__leaf_clk
rlabel metal1 s 12098 13294 12098 13294 4 clknet_2_3__leaf_clk
rlabel metal2 s 13018 959 13018 959 4 comparator_nen
rlabel metal2 s 1058 1520 1058 1520 4 dac_set[0]
rlabel metal2 s 2254 1520 2254 1520 4 dac_set[1]
rlabel metal2 s 3450 1520 3450 1520 4 dac_set[2]
rlabel metal2 s 4646 1520 4646 1520 4 dac_set[3]
rlabel metal2 s 5842 1520 5842 1520 4 dac_set[4]
rlabel metal2 s 7038 959 7038 959 4 dac_set[5]
rlabel metal2 s 8234 1520 8234 1520 4 dac_set[6]
rlabel metal2 s 9430 959 9430 959 4 dac_set[7]
rlabel metal2 s 11822 959 11822 959 4 do_calibrate
rlabel metal1 s 13013 4114 13013 4114 4 net1
rlabel metal1 s 6072 2414 6072 2414 4 net10
rlabel metal1 s 6762 4080 6762 4080 4 net11
rlabel metal1 s 8050 2414 8050 2414 4 net12
rlabel metal1 s 9798 2414 9798 2414 4 net13
rlabel metal1 s 11730 3910 11730 3910 4 net14
rlabel metal1 s 4370 13498 4370 13498 4 net15
rlabel metal3 s 3726 9044 3726 9044 4 net16
rlabel metal1 s 6210 13158 6210 13158 4 net17
rlabel metal1 s 6164 14382 6164 14382 4 net18
rlabel metal1 s 4922 14382 4922 14382 4 net19
rlabel metal4 s 12259 13804 12259 13804 4 net2
rlabel metal1 s 4094 7242 4094 7242 4 net20
rlabel metal1 s 3496 9146 3496 9146 4 net21
rlabel metal1 s 2438 14382 2438 14382 4 net22
rlabel metal1 s 1610 14348 1610 14348 4 net23
rlabel metal1 s 10672 2414 10672 2414 4 net24
rlabel metal1 s 13340 14246 13340 14246 4 net3
rlabel metal3 s 11155 13804 11155 13804 4 net4
rlabel metal1 s 12742 2414 12742 2414 4 net5
rlabel metal2 s 1610 3706 1610 3706 4 net6
rlabel metal1 s 2760 2414 2760 2414 4 net7
rlabel metal1 s 3726 2414 3726 2414 4 net8
rlabel metal1 s 4600 2414 4600 2414 4 net9
rlabel metal1 s 9200 14586 9200 14586 4 result[0]
rlabel metal1 s 8050 14586 8050 14586 4 result[1]
rlabel metal1 s 7176 14586 7176 14586 4 result[2]
rlabel metal1 s 6256 14586 6256 14586 4 result[3]
rlabel metal1 s 5152 14586 5152 14586 4 result[4]
rlabel metal1 s 4140 14586 4140 14586 4 result[5]
rlabel metal1 s 3128 14586 3128 14586 4 result[6]
rlabel metal1 s 2254 14586 2254 14586 4 result[7]
rlabel metal1 s 1242 14586 1242 14586 4 result_ready
rlabel metal1 s 13340 14382 13340 14382 4 rst
rlabel metal2 s 10626 959 10626 959 4 thresh_sel
rlabel metal3 s 10281 13668 10281 13668 4 use_ext_thresh
rlabel metal1 s 11454 14382 11454 14382 4 user_enable
flabel metal4 s 10904 2128 11304 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4904 2128 5304 14736 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7904 2128 8304 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1904 2128 2304 14736 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 14186 0 14242 800 0 FreeSans 280 90 0 0 analog_comparator_out
port 3 nsew
flabel metal2 s 12162 16589 12218 17389 0 FreeSans 280 90 0 0 calib_enable
port 4 nsew
flabel metal2 s 14186 16589 14242 17389 0 FreeSans 280 90 0 0 clk
port 5 nsew
flabel metal2 s 12990 0 13046 800 0 FreeSans 280 90 0 0 comparator_nen
port 6 nsew
flabel metal2 s 1030 0 1086 800 0 FreeSans 280 90 0 0 dac_set[0]
port 7 nsew
flabel metal2 s 2226 0 2282 800 0 FreeSans 280 90 0 0 dac_set[1]
port 8 nsew
flabel metal2 s 3422 0 3478 800 0 FreeSans 280 90 0 0 dac_set[2]
port 9 nsew
flabel metal2 s 4618 0 4674 800 0 FreeSans 280 90 0 0 dac_set[3]
port 10 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 dac_set[4]
port 11 nsew
flabel metal2 s 7010 0 7066 800 0 FreeSans 280 90 0 0 dac_set[5]
port 12 nsew
flabel metal2 s 8206 0 8262 800 0 FreeSans 280 90 0 0 dac_set[6]
port 13 nsew
flabel metal2 s 9402 0 9458 800 0 FreeSans 280 90 0 0 dac_set[7]
port 14 nsew
flabel metal2 s 11794 0 11850 800 0 FreeSans 280 90 0 0 do_calibrate
port 15 nsew
flabel metal2 s 9126 16589 9182 17389 0 FreeSans 280 90 0 0 result[0]
port 16 nsew
flabel metal2 s 8114 16589 8170 17389 0 FreeSans 280 90 0 0 result[1]
port 17 nsew
flabel metal2 s 7102 16589 7158 17389 0 FreeSans 280 90 0 0 result[2]
port 18 nsew
flabel metal2 s 6090 16589 6146 17389 0 FreeSans 280 90 0 0 result[3]
port 19 nsew
flabel metal2 s 5078 16589 5134 17389 0 FreeSans 280 90 0 0 result[4]
port 20 nsew
flabel metal2 s 4066 16589 4122 17389 0 FreeSans 280 90 0 0 result[5]
port 21 nsew
flabel metal2 s 3054 16589 3110 17389 0 FreeSans 280 90 0 0 result[6]
port 22 nsew
flabel metal2 s 2042 16589 2098 17389 0 FreeSans 280 90 0 0 result[7]
port 23 nsew
flabel metal2 s 1030 16589 1086 17389 0 FreeSans 280 90 0 0 result_ready
port 24 nsew
flabel metal2 s 13174 16589 13230 17389 0 FreeSans 280 90 0 0 rst
port 25 nsew
flabel metal2 s 10598 0 10654 800 0 FreeSans 280 90 0 0 thresh_sel
port 26 nsew
flabel metal2 s 10138 16589 10194 17389 0 FreeSans 280 90 0 0 use_ext_thresh
port 27 nsew
flabel metal2 s 11150 16589 11206 17389 0 FreeSans 280 90 0 0 user_enable
port 28 nsew
<< properties >>
string FIXED_BBOX 0 0 15245 17389
string GDS_END 1023298
string GDS_FILE wowa_digital.gds
string GDS_START 374716
<< end >>
