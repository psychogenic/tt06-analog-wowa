* NGSPICE file created from calibrated_comparator_parax.ext - technology: sky130A

.subckt calibrated_comparator_parax INPUT VCC THRESHV VSS CALIB RESULT EN_N
X0 x3.OUT.t2 x3.SEL_N.t2 INPUT.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X1 x1.inhigh.t0 THRESHV.t2 x1.G1 VCC.t0 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=2.32 ps=17.03111 w=8 l=2
**devattr s=92800,3316 d=92800,3316
X2 x2.OUT.t2 VSS.t9 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 THRESHV.t1 x3.SEL_N.t3 x3.OUT.t3 VCC sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X4 VCC.t6 EN_N.t0 x1.p2p VCC.t5 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=8
**devattr s=11600,516 d=11600,516
X5 x1.G2 x3.OUT.t4 x1.inhigh.t1 VCC.t9 sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=0 ps=0 w=8 l=2
**devattr s=92800,3316 d=92800,3316
X6 x2.x2.Z VSS.t7 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 x1.pg2g x1.G1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=4
**devattr s=23200,916 d=23200,916
X8 VSS.t5 EN_N.t1 RESULT.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X9 x1.mirhigh.t1 x1.pg2g.t2 RESULT.t3 VCC.t10 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=4
**devattr s=46400,1716 d=46400,1716
X10 x3.OUT.t1 CALIB.t0 INPUT.t0 VCC sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X11 VSS.t16 x1.G2 RESULT.t1 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=4
**devattr s=23200,916 d=23200,916
X12 x1.pg2g.t1 x1.pg2g.t0 x1.mirhigh.t2 VCC.t7 sky130_fd_pr__pfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=4 l=4
**devattr s=46400,1716 d=46400,1716
X13 x2.x2.GP CALIB.t1 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X14 x2.OUT.t2 VSS.t8 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X15 x1.n2n VCC.t15 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=8
**devattr s=5800,316 d=5800,316
X16 x3.SEL_N.t1 CALIB.t2 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=11600,516 d=11600,516
X17 VSS.t1 x1.G1 x1.G1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0.58 ps=4.928 w=2 l=4
**devattr s=23200,916 d=23200,916
X18 x2.OUT.t0 CALIB.t3 RESULT.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X19 x1.inhigh.t2 EN_N.t2 VCC.t14 VCC.t13 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=8
**devattr s=23200,916 d=23200,916
X20 VCC CALIB.t4 x2.x2.GP VCC sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=13.45 as=0.58 ps=4.58 w=2 l=0.35
**devattr s=23200,916 d=23200,916
X21 VCC.t12 EN_N.t3 x1.mirhigh.t0 VCC.t11 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=0.15
**devattr s=58000,2116 d=58000,2116
X22 VCC CALIB.t5 x3.SEL_N.t0 VCC sky130_fd_pr__pfet_01v8_lvt ad=1.74 pd=13.45 as=0 ps=0 w=2 l=0.35
**devattr s=23200,916 d=23200,916
X23 x1.G1 x2.OUT.t3 x1.p2p VCC.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.128889 as=0.29 ps=2.58 w=1 l=1
**devattr s=11600,516 d=11600,516
X24 x1.G1 x2.OUT.t4 x1.n2n VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.232 as=0.145 ps=1.58 w=0.5 l=1
**devattr s=5800,316 d=5800,316
X25 x1.G2 x1.G2 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0 ps=0 w=2 l=4
**devattr s=23200,916 d=23200,916
X26 THRESHV.t0 CALIB.t6 x3.OUT.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X27 x2.OUT.t1 x2.x2.GP RESULT.t4 VCC sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.2
**devattr s=23200,916 d=23200,916
X28 x2.x2.Z VSS.t6 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
R0 x3.x2.GP x3.SEL_N.t3 239.171
R1 x3.x3.GN x3.SEL_N.t2 233.901
R2 x3.x2.GP x3.SEL_N.t0 113.802
R3 x3.x2.GP x3.SEL_N.t1 83.8505
R4 x3.x2.GP x3.x3.GN 6.46588
R5 INPUT.n1 INPUT.t0 113.761
R6 INPUT INPUT.t1 41.5734
R7 INPUT.n2 INPUT 0.724136
R8 INPUT INPUT.n1 0.272792
R9 INPUT.n1 INPUT.n0 0.0970909
R10 INPUT.n0 INPUT 0.08175
R11 INPUT.n2 INPUT 0.06925
R12 INPUT INPUT.n2 0.063
R13 INPUT.n0 INPUT 0.0573182
R14 x3.OUT x3.OUT.t1 113.803
R15 x3.OUT x3.OUT.t3 113.796
R16 x3.OUT x3.OUT.t4 68.4234
R17 x3.OUT x3.OUT.t0 41.6342
R18 x3.OUT x3.OUT.t2 41.507
R19 x3.OUT x3.OUT.n0 7.4523
R20 x3.OUT.n0 x3.OUT 2.78298
R21 x3.OUT.n0 x3.OUT 1.90525
R22 x3.OUT.n0 x3.OUT 1.89141
R23 VSS.n174 VSS.n173 88402
R24 VSS.n65 VSS.n10 54813.6
R25 VSS.n223 VSS.n10 23373.5
R26 VSS.n173 VSS.n172 20661.8
R27 VSS.n167 VSS.n166 20589.7
R28 VSS.n223 VSS.n9 20389.3
R29 VSS.n166 VSS.n103 19594.2
R30 VSS.n173 VSS.n170 16402.4
R31 VSS.n170 VSS.n75 15575.6
R32 VSS.n101 VSS.n100 15459.7
R33 VSS.n170 VSS.n169 14979.4
R34 VSS.n169 VSS.n168 14273.2
R35 VSS.n100 VSS.n76 11532
R36 VSS.n166 VSS.n165 10139.7
R37 VSS.n102 VSS.n101 8515.32
R38 VSS.n171 VSS.n9 8485.71
R39 VSS.n101 VSS.n75 8450.84
R40 VSS.n100 VSS.n99 7837.4
R41 VSS.n165 VSS.n102 7359.64
R42 VSS.n167 VSS.n102 7196.9
R43 VSS.n89 VSS.n77 6564.74
R44 VSS.n98 VSS.n77 6564.74
R45 VSS.n89 VSS.n78 6564.74
R46 VSS.n98 VSS.n78 6564.74
R47 VSS.n211 VSS.n22 5178.05
R48 VSS.n148 VSS.n56 5116.21
R49 VSS.n189 VSS.n56 5116.21
R50 VSS.n148 VSS.n57 5116.21
R51 VSS.n189 VSS.n57 5116.21
R52 VSS.n179 VSS.n63 5116.21
R53 VSS.n179 VSS.n64 5116.21
R54 VSS.n180 VSS.n64 5116.21
R55 VSS.n180 VSS.n63 5116.21
R56 VSS.n129 VSS.n110 5116.21
R57 VSS.n150 VSS.n110 5116.21
R58 VSS.n150 VSS.n111 5116.21
R59 VSS.n129 VSS.n111 5116.21
R60 VSS.n175 VSS.n5 5116.21
R61 VSS.n225 VSS.n5 5116.21
R62 VSS.n175 VSS.n6 5116.21
R63 VSS.n225 VSS.n6 5116.21
R64 VSS.n164 VSS.n163 4543.31
R65 VSS.n165 VSS.n164 3590.61
R66 VSS.n99 VSS.n22 3277.63
R67 VSS.n33 VSS.n29 2914.44
R68 VSS.n41 VSS.n29 2914.44
R69 VSS.n41 VSS.n30 2914.44
R70 VSS.n33 VSS.n30 2914.44
R71 VSS.n162 VSS.n105 2914.44
R72 VSS.n155 VSS.n105 2914.44
R73 VSS.n162 VSS.n106 2914.44
R74 VSS.n155 VSS.n106 2914.44
R75 VSS.n210 VSS.n18 2914.44
R76 VSS.n210 VSS.n19 2914.44
R77 VSS.n213 VSS.n19 2914.44
R78 VSS.n213 VSS.n18 2914.44
R79 VSS.n192 VSS.n191 2837.13
R80 VSS.n21 VSS.n20 2519.66
R81 VSS.n92 VSS.n83 2508.85
R82 VSS.n92 VSS.n84 2508.85
R83 VSS.n93 VSS.n83 2508.85
R84 VSS.n93 VSS.n84 2508.85
R85 VSS.n169 VSS.n167 2472.45
R86 VSS.n221 VSS.n11 2306.06
R87 VSS.n38 VSS.n11 2306.06
R88 VSS.n221 VSS.n12 2306.06
R89 VSS.n38 VSS.n12 2306.06
R90 VSS.n120 VSS.n119 2306.06
R91 VSS.n132 VSS.n119 2306.06
R92 VSS.n128 VSS.n120 2306.06
R93 VSS.n132 VSS.n128 2306.06
R94 VSS.n194 VSS.n52 2306.06
R95 VSS.n194 VSS.n53 2306.06
R96 VSS.n195 VSS.n52 2306.06
R97 VSS.n195 VSS.n53 2306.06
R98 VSS.n22 VSS.n21 2129.58
R99 VSS.n191 VSS.n10 2068.85
R100 VSS.n174 VSS.t0 1874.46
R101 VSS.n90 VSS.n89 1872.69
R102 VSS.n90 VSS.t11 1789.83
R103 VSS.n153 VSS.n54 1658.64
R104 VSS.n85 VSS.n75 1577.45
R105 VSS.n164 VSS.n104 1382.33
R106 VSS.n153 VSS.n152 1314.03
R107 VSS.t20 VSS.n54 1285
R108 VSS.t20 VSS.n192 1285
R109 VSS.t23 VSS.n85 1137.45
R110 VSS.n154 VSS.n153 996.365
R111 VSS.n90 VSS.n76 856.596
R112 VSS.n35 VSS.n34 761.481
R113 VSS.n39 VSS.n20 706.557
R114 VSS.n225 VSS.n224 696.282
R115 VSS.t13 VSS.n66 678.75
R116 VSS.n163 VSS.t17 592.727
R117 VSS.n154 VSS.t17 592.727
R118 VSS.n212 VSS.n20 553.96
R119 VSS.n131 VSS.n130 514.71
R120 VSS.n130 VSS.t15 502.255
R121 VSS.n147 VSS.t2 502.144
R122 VSS.n178 VSS.n67 451.89
R123 VSS.n40 VSS.t18 450.954
R124 VSS.n223 VSS.n7 441.522
R125 VSS.n152 VSS.n151 435.562
R126 VSS.n88 VSS.n79 426.541
R127 VSS.n176 VSS.n74 426.505
R128 VSS.n212 VSS.t22 389.784
R129 VSS.t22 VSS.n211 389.784
R130 VSS.n97 VSS.n79 359.279
R131 VSS.n188 VSS.n58 322.786
R132 VSS.n223 VSS.n222 312.2
R133 VSS.n191 VSS.t2 298.697
R134 VSS.n224 VSS.t0 292.769
R135 VSS.n53 VSS.n51 292.5
R136 VSS.n192 VSS.n53 292.5
R137 VSS.n52 VSS.n50 292.5
R138 VSS.n54 VSS.n52 292.5
R139 VSS.n23 VSS.n18 292.5
R140 VSS.t22 VSS.n18 292.5
R141 VSS.n24 VSS.n19 292.5
R142 VSS.t22 VSS.n19 292.5
R143 VSS.n128 VSS.n127 292.5
R144 VSS.t4 VSS.n128 292.5
R145 VSS.n123 VSS.n119 292.5
R146 VSS.t4 VSS.n119 292.5
R147 VSS.n108 VSS.n106 292.5
R148 VSS.n106 VSS.t17 292.5
R149 VSS.n107 VSS.n105 292.5
R150 VSS.n105 VSS.t17 292.5
R151 VSS.n34 VSS.n33 292.5
R152 VSS.n33 VSS.n9 292.5
R153 VSS.n42 VSS.n41 292.5
R154 VSS.n41 VSS.n40 292.5
R155 VSS.n38 VSS.n37 292.5
R156 VSS.n39 VSS.n38 292.5
R157 VSS.n221 VSS.n220 292.5
R158 VSS.n222 VSS.n221 292.5
R159 VSS.t23 VSS.n90 280.851
R160 VSS.n222 VSS.t10 268.382
R161 VSS.n183 VSS.n62 258.839
R162 VSS.n178 VSS.n177 249.601
R163 VSS.n177 VSS.n176 249.601
R164 VSS.n226 VSS.n4 244.138
R165 VSS.t11 VSS.n22 238.644
R166 VSS.n96 VSS.t12 229.185
R167 VSS.n122 VSS.n121 217.103
R168 VSS.n224 VSS.n223 206.661
R169 VSS.n191 VSS.n190 203.447
R170 VSS.t18 VSS.t10 200.831
R171 VSS.n121 VSS.n112 198.024
R172 VSS.n112 VSS.n58 198.024
R173 VSS.n190 VSS.n55 197.899
R174 VSS.n156 VSS.n107 189.365
R175 VSS.n161 VSS.n107 189.365
R176 VSS.t13 VSS.n65 183.857
R177 VSS.n157 VSS.n156 181.929
R178 VSS.n151 VSS.n103 177.554
R179 VSS.t4 VSS.n104 171.571
R180 VSS.n131 VSS.t4 171.571
R181 VSS.n91 VSS.n82 163.012
R182 VSS.n91 VSS.n81 163.012
R183 VSS.n94 VSS.n82 158.72
R184 VSS.n95 VSS.n81 156.988
R185 VSS.n168 VSS.n65 151.661
R186 VSS.n193 VSS.n51 149.835
R187 VSS.n193 VSS.n50 149.835
R188 VSS.n220 VSS.n13 149.835
R189 VSS.n147 VSS.n103 149.811
R190 VSS.n98 VSS.n97 146.25
R191 VSS.n99 VSS.n98 146.25
R192 VSS.n89 VSS.n88 146.25
R193 VSS.n84 VSS.n82 146.25
R194 VSS.n84 VSS.n76 146.25
R195 VSS.n83 VSS.n81 146.25
R196 VSS.n85 VSS.n83 146.25
R197 VSS.n67 VSS.n62 140.8
R198 VSS.n37 VSS.n13 129.781
R199 VSS.n196 VSS.n51 126.947
R200 VSS.n74 VSS.n4 126.721
R201 VSS.n197 VSS.n50 124.462
R202 VSS.n194 VSS.n193 117.001
R203 VSS.t20 VSS.n194 117.001
R204 VSS.n196 VSS.n195 117.001
R205 VSS.n195 VSS.t20 117.001
R206 VSS.n133 VSS.n132 117.001
R207 VSS.n132 VSS.n131 117.001
R208 VSS.n125 VSS.n120 117.001
R209 VSS.n120 VSS.n104 117.001
R210 VSS.n14 VSS.n12 117.001
R211 VSS.t18 VSS.n12 117.001
R212 VSS.n13 VSS.n11 117.001
R213 VSS.t18 VSS.n11 117.001
R214 VSS.n92 VSS.n91 117.001
R215 VSS.t23 VSS.n92 117.001
R216 VSS.n94 VSS.n93 117.001
R217 VSS.n93 VSS.t23 117.001
R218 VSS.n161 VSS.n160 91.8593
R219 VSS.n115 VSS.t5 86.7387
R220 VSS.n160 VSS.n108 85.9864
R221 VSS.n199 VSS.t21 83.7422
R222 VSS.n218 VSS.t19 83.7278
R223 VSS.n29 VSS.n16 77.0112
R224 VSS.n209 VSS.n23 76.5461
R225 VSS.n34 VSS.n32 76.3348
R226 VSS.n187 VSS.n59 76.1229
R227 VSS.n177 VSS.n68 75.9791
R228 VSS.n73 VSS.n5 75.6884
R229 VSS.n210 VSS.n209 73.1255
R230 VSS.n211 VSS.n210 73.1255
R231 VSS.n214 VSS.n213 73.1255
R232 VSS.n213 VSS.n212 73.1255
R233 VSS.n129 VSS.n118 73.1255
R234 VSS.n130 VSS.n129 73.1255
R235 VSS.n156 VSS.n155 73.1255
R236 VSS.n155 VSS.n154 73.1255
R237 VSS.n162 VSS.n161 73.1255
R238 VSS.n163 VSS.n162 73.1255
R239 VSS.n67 VSS.n63 73.1255
R240 VSS.n63 VSS.n55 73.1255
R241 VSS.n150 VSS.n149 73.1255
R242 VSS.n151 VSS.n150 73.1255
R243 VSS.n189 VSS.n188 73.1255
R244 VSS.n190 VSS.n189 73.1255
R245 VSS.n149 VSS.n148 73.1255
R246 VSS.n148 VSS.n147 73.1255
R247 VSS.n68 VSS.n64 73.1255
R248 VSS.n66 VSS.n64 73.1255
R249 VSS.n8 VSS.n5 73.1255
R250 VSS.n32 VSS.n30 73.1255
R251 VSS.n30 VSS.t10 73.1255
R252 VSS.n29 VSS.t10 73.1255
R253 VSS.n74 VSS.n6 73.1255
R254 VSS.n7 VSS.n6 73.1255
R255 VSS.n88 VSS.n87 71.5299
R256 VSS.n152 VSS.t15 66.5831
R257 VSS.n31 VSS.n23 65.1299
R258 VSS.n172 VSS.n171 65.0005
R259 VSS.n124 VSS.n123 54.9719
R260 VSS.n220 VSS.n219 53.4638
R261 VSS.n87 VSS.n4 53.3135
R262 VSS.n171 VSS.n8 50.0005
R263 VSS.n226 VSS.n225 41.7862
R264 VSS.n176 VSS.n175 41.7862
R265 VSS.n175 VSS.n174 41.7862
R266 VSS.n143 VSS.n111 41.7862
R267 VSS.n111 VSS.t15 41.7862
R268 VSS.n121 VSS.n110 41.7862
R269 VSS.n110 VSS.t15 41.7862
R270 VSS.n145 VSS.n57 41.7862
R271 VSS.n57 VSS.t2 41.7862
R272 VSS.n58 VSS.n56 41.7862
R273 VSS.n56 VSS.t2 41.7862
R274 VSS.n181 VSS.n180 41.7862
R275 VSS.n180 VSS.t13 41.7862
R276 VSS.n179 VSS.n178 41.7862
R277 VSS.t13 VSS.n179 41.7862
R278 VSS.n114 VSS.t16 41.7156
R279 VSS.n69 VSS.t14 41.4575
R280 VSS.n71 VSS.t1 41.4563
R281 VSS.n186 VSS.t3 41.4498
R282 VSS.n134 VSS.n117 39.1319
R283 VSS.n134 VSS.n133 38.7101
R284 VSS.n126 VSS.n125 37.7441
R285 VSS.n72 VSS.n3 34.0553
R286 VSS.n127 VSS.n126 32.9148
R287 VSS.n168 VSS.n55 30.5175
R288 VSS.n177 VSS.n73 26.3819
R289 VSS.n209 VSS.n208 24.5021
R290 VSS.n86 VSS.n78 23.4005
R291 VSS.t11 VSS.n78 23.4005
R292 VSS.n79 VSS.n77 23.4005
R293 VSS.t11 VSS.n77 23.4005
R294 VSS.n188 VSS.n187 21.7605
R295 VSS.n223 VSS.n8 20.0005
R296 VSS.n124 VSS.n116 19.81
R297 VSS.n40 VSS.n39 18.2578
R298 VSS.n181 VSS.n3 16.6656
R299 VSS.n123 VSS.n122 16.4078
R300 VSS.n227 VSS.n3 16.3973
R301 VSS.n172 VSS.n66 15.0005
R302 VSS.n32 VSS.n26 13.4459
R303 VSS.n149 VSS.n112 11.5469
R304 VSS.n149 VSS.n146 11.217
R305 VSS.n37 VSS.n36 10.4904
R306 VSS.n183 VSS.n182 10.4191
R307 VSS.n97 VSS.n80 10.2128
R308 VSS.n125 VSS.n124 9.84665
R309 VSS.n45 VSS.n44 9.39185
R310 VSS.n135 VSS.n116 9.37653
R311 VSS.n49 VSS.n26 9.363
R312 VSS.n28 VSS.n24 9.3445
R313 VSS.n160 VSS.n159 9.3005
R314 VSS.n97 VSS.n96 9.3005
R315 VSS.n80 VSS.n1 7.99658
R316 VSS.n87 VSS.n86 7.45136
R317 VSS.n126 VSS.n116 7.13193
R318 VSS.n96 VSS.n95 6.74718
R319 VSS.n122 VSS.n118 6.4257
R320 VSS.n146 VSS.n143 6.18574
R321 VSS.n146 VSS.n145 6.18574
R322 VSS.n36 VSS.n31 5.33383
R323 VSS.n134 VSS.n113 4.90573
R324 VSS.n43 VSS.n26 4.84084
R325 VSS.n144 VSS.n59 4.59111
R326 VSS.n36 VSS.n35 4.44494
R327 VSS.n72 VSS.n68 4.36414
R328 VSS.n21 VSS.n7 3.80673
R329 VSS.n35 VSS.n16 3.68304
R330 VSS.n36 VSS.n14 3.37828
R331 VSS.n143 VSS.n142 3.29929
R332 VSS.n72 VSS.n69 3.1005
R333 VSS.n72 VSS.n71 3.1005
R334 VSS.n44 VSS.n43 3.04897
R335 VSS.n31 VSS.n16 3.03114
R336 VSS.n214 VSS.n17 2.76373
R337 VSS.n208 VSS.n207 2.3255
R338 VSS.n17 VSS.n15 2.3255
R339 VSS.n158 VSS.n157 2.3255
R340 VSS.n117 VSS.n115 1.89317
R341 VSS.n215 VSS.n16 1.87237
R342 VSS.n219 VSS.n218 1.86348
R343 VSS.n198 VSS.n197 1.8605
R344 VSS.n187 VSS.n186 1.8605
R345 VSS.n114 VSS.n113 1.8605
R346 VSS.n62 VSS.n59 1.85321
R347 VSS.n44 VSS.n42 1.67627
R348 VSS.n135 VSS.n134 1.66708
R349 VSS.n73 VSS.n72 1.46981
R350 VSS.n216 VSS.n215 1.32907
R351 VSS.n197 VSS.n196 1.2805
R352 VSS.n95 VSS.n94 1.2805
R353 VSS.n203 VSS 1.2505
R354 VSS.n231 VSS 1.2505
R355 VSS.n137 VSS.t8 1.21428
R356 VSS.n138 VSS.t6 1.21428
R357 VSS.n186 VSS.n185 1.06892
R358 VSS.n138 VSS.n137 1.04896
R359 VSS.n133 VSS.n118 1.00837
R360 VSS.n215 VSS.n214 0.981001
R361 VSS.n201 VSS 0.976194
R362 VSS.n46 VSS.n28 0.939674
R363 VSS.n159 VSS.t6 0.909702
R364 VSS.n182 VSS.n61 0.845955
R365 VSS.n228 VSS.n227 0.845955
R366 VSS.n144 VSS.n60 0.592183
R367 VSS.n229 VSS.n1 0.529939
R368 VSS.n140 VSS.n60 0.520386
R369 VSS.n142 VSS.n141 0.517167
R370 VSS.n136 VSS.n135 0.517167
R371 VSS.n80 VSS.n0 0.517167
R372 VSS.n139 VSS.t7 0.473714
R373 VSS.n229 VSS.n228 0.462148
R374 VSS.n204 VSS.n202 0.407111
R375 VSS.n96 VSS.n0 0.405672
R376 VSS.n204 VSS.n203 0.367895
R377 VSS.n43 VSS.n28 0.339219
R378 VSS.n157 VSS.n108 0.3205
R379 VSS VSS.n109 0.315747
R380 VSS.n182 VSS.n181 0.268407
R381 VSS.n227 VSS.n226 0.268407
R382 VSS.n217 VSS.n216 0.263801
R383 VSS VSS.n229 0.236295
R384 VSS.n140 VSS.n139 0.21925
R385 VSS.n218 VSS.n217 0.197673
R386 VSS.n230 VSS.n0 0.194466
R387 VSS.n86 VSS.n1 0.188758
R388 VSS.n127 VSS.n117 0.183357
R389 VSS.n201 VSS.n49 0.172797
R390 VSS.n61 VSS.n2 0.172375
R391 VSS.n228 VSS.n2 0.166693
R392 VSS.n137 VSS.t9 0.165823
R393 VSS.t7 VSS.n138 0.165823
R394 VSS.n141 VSS.n114 0.163852
R395 VSS.n48 VSS.n27 0.15675
R396 VSS.n205 VSS 0.154346
R397 VSS.n202 VSS.n25 0.152527
R398 VSS.n136 VSS.n115 0.151068
R399 VSS.n70 VSS.n2 0.146333
R400 VSS.n185 VSS.n60 0.141125
R401 VSS.n139 VSS.n136 0.136864
R402 VSS.n141 VSS.n140 0.128341
R403 VSS.n205 VSS 0.1255
R404 VSS.n185 VSS.n184 0.122659
R405 VSS.n200 VSS 0.113
R406 VSS.n202 VSS.n201 0.108139
R407 VSS.n184 VSS.n61 0.0999318
R408 VSS.n231 VSS.n230 0.0999318
R409 VSS.n47 VSS.n46 0.0957944
R410 VSS.n216 VSS.n15 0.0954519
R411 VSS.n200 VSS.n199 0.0934487
R412 VSS.n198 VSS 0.088641
R413 VSS.n49 VSS.n48 0.0861481
R414 VSS VSS.n204 0.0835761
R415 VSS.n145 VSS.n144 0.0729516
R416 VSS.n159 VSS.n158 0.0684987
R417 VSS.n208 VSS.n24 0.0645
R418 VSS.n207 VSS.n25 0.063
R419 VSS.n230 VSS 0.0558977
R420 VSS.n45 VSS.n25 0.0540714
R421 VSS.n158 VSS 0.0518393
R422 VSS.n219 VSS.n14 0.0512937
R423 VSS.n217 VSS 0.047375
R424 VSS.n184 VSS.n183 0.047
R425 VSS.n142 VSS.n113 0.043453
R426 VSS.n47 VSS 0.0411786
R427 VSS.n109 VSS 0.0402727
R428 VSS VSS.n200 0.0325513
R429 VSS.n206 VSS 0.03175
R430 VSS.n70 VSS.n69 0.03175
R431 VSS.n71 VSS.n70 0.03175
R432 VSS.n109 VSS 0.0229359
R433 VSS.n207 VSS.n206 0.0205893
R434 VSS.n27 VSS.n15 0.0205893
R435 VSS.n46 VSS.n45 0.0192927
R436 VSS.n27 VSS 0.0183571
R437 VSS.n42 VSS.n17 0.0183273
R438 VSS.n48 VSS.n47 0.0152857
R439 VSS.n206 VSS.n205 0.0101154
R440 VSS.n203 VSS 0.00387838
R441 VSS VSS.n231 0.00334091
R442 VSS.n199 VSS.n198 0.00210256
R443 THRESHV.n1 THRESHV.t1 113.788
R444 THRESHV.n4 THRESHV.t2 68.4093
R445 THRESHV THRESHV.t0 41.5734
R446 THRESHV.n5 THRESHV.n4 8.95852
R447 THRESHV.n2 THRESHV.n1 8.3611
R448 THRESHV.n5 THRESHV 0.226603
R449 THRESHV THRESHV.n5 0.142044
R450 THRESHV.n3 THRESHV 0.1255
R451 THRESHV.n0 THRESHV 0.0966538
R452 THRESHV.n2 THRESHV 0.0609346
R453 THRESHV.n0 THRESHV 0.0573182
R454 THRESHV.n4 THRESHV 0.0236642
R455 THRESHV.n1 THRESHV.n0 0.0175455
R456 THRESHV THRESHV.n3 0.0170441
R457 THRESHV.n3 THRESHV.n2 0.0126344
R458 x1.inhigh x1.inhigh.t2 115.745
R459 x1.inhigh x1.inhigh.t1 31.1787
R460 x1.inhigh x1.inhigh.t0 29.4286
R461 VCC.n88 VCC.n87 4560
R462 VCC.n85 VCC.n83 4560
R463 VCC.n73 VCC.n70 4560
R464 VCC.n76 VCC.n69 4560
R465 VCC.n34 VCC.n32 4560
R466 VCC.n37 VCC.n36 4560
R467 VCC.n101 VCC.n15 4207.06
R468 VCC.n98 VCC.n16 4207.06
R469 VCC.n49 VCC.n43 3854.12
R470 VCC.n47 VCC.n46 3854.12
R471 VCC.n26 VCC.n25 3854.12
R472 VCC.n23 VCC.n21 3854.12
R473 VCC.n62 VCC.n56 2848.24
R474 VCC.n60 VCC.n59 2848.24
R475 VCC.n9 VCC.n8 1736.47
R476 VCC.n6 VCC.n4 1736.47
R477 VCC.n99 VCC.n15 1068.61
R478 VCC.n100 VCC.n16 1068.61
R479 VCC.n59 VCC.n58 1018.62
R480 VCC.n62 VCC.n61 1018.62
R481 VCC.n74 VCC.n69 879.971
R482 VCC.n75 VCC.n70 879.971
R483 VCC.n84 VCC.n80 486.401
R484 VCC.n84 VCC.n81 486.401
R485 VCC.n89 VCC.n81 486.401
R486 VCC.n77 VCC.n68 486.401
R487 VCC.n33 VCC.n29 486.401
R488 VCC.n33 VCC.n30 486.401
R489 VCC.n38 VCC.n30 486.401
R490 VCC.n78 VCC.n77 468.406
R491 VCC.n102 VCC.n14 443.728
R492 VCC.n103 VCC.n102 436.236
R493 VCC.n50 VCC.n42 411.106
R494 VCC.n44 VCC.n42 411.106
R495 VCC.n22 VCC.n18 411.106
R496 VCC.n22 VCC.n19 411.106
R497 VCC.n44 VCC.n41 387.128
R498 VCC.n46 VCC.n45 385.567
R499 VCC.n49 VCC.n48 385.567
R500 VCC.n26 VCC.n20 385.567
R501 VCC.n24 VCC.n23 385.567
R502 VCC.n51 VCC.n50 384.087
R503 VCC.n27 VCC.n19 354.171
R504 VCC.n72 VCC.n67 349.312
R505 VCC.n71 VCC.n68 333.82
R506 VCC.n28 VCC.n18 321.255
R507 VCC.n9 VCC.n3 314.781
R508 VCC.n7 VCC.n6 314.781
R509 VCC.n63 VCC.n55 303.812
R510 VCC.n57 VCC.n55 303.812
R511 VCC.n97 VCC.n17 285.354
R512 VCC.n96 VCC.n13 272.99
R513 VCC.n90 VCC.n89 265.865
R514 VCC.n39 VCC.n29 249.901
R515 VCC.n91 VCC.t6 228.284
R516 VCC.n57 VCC.n54 215.555
R517 VCC.n64 VCC.n63 213.397
R518 VCC.n90 VCC.n80 186.805
R519 VCC.n39 VCC.n38 185.901
R520 VCC.n5 VCC.n1 185.225
R521 VCC.n5 VCC.n2 185.225
R522 VCC.n10 VCC.n2 162.456
R523 VCC.n88 VCC.n82 160.32
R524 VCC.n86 VCC.n85 160.32
R525 VCC.n35 VCC.n34 160.32
R526 VCC.n37 VCC.n31 160.32
R527 VCC.n11 VCC.n1 159.474
R528 VCC.n79 VCC.t14 113.716
R529 VCC.n63 VCC.n62 92.5005
R530 VCC.n59 VCC.n57 92.5005
R531 VCC.n53 VCC.t12 48.1635
R532 VCC.n4 VCC.n1 37.0005
R533 VCC.n8 VCC.n2 37.0005
R534 VCC.n16 VCC.n14 30.8338
R535 VCC.n15 VCC.n13 30.8338
R536 VCC.n6 VCC.n5 30.8338
R537 VCC.n10 VCC.n9 30.8338
R538 VCC.n4 VCC.n3 29.6618
R539 VCC.n8 VCC.n7 29.6618
R540 VCC.n83 VCC.n80 23.1255
R541 VCC.n87 VCC.n81 23.1255
R542 VCC.n70 VCC.n67 23.1255
R543 VCC.n69 VCC.n68 23.1255
R544 VCC.n32 VCC.n29 23.1255
R545 VCC.n36 VCC.n30 23.1255
R546 VCC.n83 VCC.n82 22.2004
R547 VCC.n87 VCC.n86 22.2004
R548 VCC.n32 VCC.n31 22.2004
R549 VCC.n36 VCC.n35 22.2004
R550 VCC.n50 VCC.n49 13.2148
R551 VCC.n47 VCC.n42 13.2148
R552 VCC.n46 VCC.n44 13.2148
R553 VCC.n43 VCC.n41 13.2148
R554 VCC.n21 VCC.n18 13.2148
R555 VCC.n23 VCC.n22 13.2148
R556 VCC.n25 VCC.n19 13.2148
R557 VCC.n27 VCC.n26 13.2148
R558 VCC.n28 VCC.n27 13.0138
R559 VCC.n45 VCC.n43 11.8527
R560 VCC.n48 VCC.n47 11.8527
R561 VCC.n21 VCC.n20 11.8527
R562 VCC.n25 VCC.n24 11.8527
R563 VCC.n60 VCC.n55 10.8829
R564 VCC.n56 VCC.n54 10.8829
R565 VCC.n72 VCC.n71 9.08437
R566 VCC.n12 VCC.t15 8.96809
R567 VCC.n77 VCC.n76 7.4005
R568 VCC.n73 VCC.n72 7.4005
R569 VCC.n98 VCC.n97 7.4005
R570 VCC.n102 VCC.n101 7.4005
R571 VCC.n85 VCC.n84 7.11588
R572 VCC.n89 VCC.n88 7.11588
R573 VCC.n34 VCC.n33 7.11588
R574 VCC.n38 VCC.n37 7.11588
R575 VCC.n58 VCC.n56 6.96486
R576 VCC.n61 VCC.n60 6.96486
R577 VCC.n7 VCC.t8 6.70818
R578 VCC.t8 VCC.n3 6.70818
R579 VCC.n74 VCC.n73 5.9633
R580 VCC.n76 VCC.n75 5.9633
R581 VCC.n99 VCC.n98 5.51167
R582 VCC.n101 VCC.n100 5.51167
R583 VCC.n95 VCC.n94 4.96483
R584 VCC.n78 VCC.n67 4.8645
R585 VCC.n61 VCC.t11 3.89288
R586 VCC.n58 VCC.t11 3.89288
R587 VCC.n52 VCC.n40 3.72362
R588 VCC.n79 VCC.n78 3.1005
R589 VCC.n91 VCC.n17 3.1005
R590 VCC.n97 VCC.n96 2.84494
R591 VCC.n92 VCC.n90 2.6261
R592 VCC.n52 VCC.n51 1.9301
R593 VCC.n17 VCC.n14 1.9205
R594 VCC.n100 VCC.t5 1.88064
R595 VCC.t5 VCC.n99 1.88064
R596 VCC.n12 VCC.n11 1.8605
R597 VCC.n104 VCC.n103 1.8605
R598 VCC.n40 VCC.n39 1.663
R599 VCC.n11 VCC.n10 1.5365
R600 VCC.n51 VCC.n41 1.47742
R601 VCC.n75 VCC.t13 1.42902
R602 VCC.t13 VCC.n74 1.42902
R603 VCC.n48 VCC.t10 1.32296
R604 VCC.n45 VCC.t10 1.32296
R605 VCC.n24 VCC.t7 1.32296
R606 VCC.t7 VCC.n20 1.32296
R607 VCC.n103 VCC.n13 1.2805
R608 VCC.n64 VCC.n54 0.853833
R609 VCC.n40 VCC.n28 0.846486
R610 VCC.n86 VCC.t0 0.814017
R611 VCC.t0 VCC.n82 0.814017
R612 VCC.t9 VCC.n31 0.814017
R613 VCC.n35 VCC.t9 0.814017
R614 VCC.n65 VCC.n64 0.6205
R615 VCC.n66 VCC.n65 0.510369
R616 VCC.n53 VCC.n52 0.490955
R617 VCC.n104 VCC.n12 0.429597
R618 VCC.n71 VCC.n66 0.423227
R619 VCC.n96 VCC.n95 0.423227
R620 VCC.n94 VCC.n66 0.321523
R621 VCC.n0 VCC 0.303385
R622 VCC.n93 VCC.n92 0.280262
R623 VCC.n94 VCC.n93 0.224184
R624 VCC VCC.n104 0.169416
R625 VCC.n92 VCC.n91 0.140381
R626 VCC VCC.n0 0.0946265
R627 VCC.n93 VCC.n79 0.0268158
R628 VCC.n95 VCC.n0 0.0178193
R629 VCC.n65 VCC.n53 0.00130906
R630 x2.x2.Z x2.OUT.t1 113.781
R631 x1.ADJ x2.OUT.t3 60.56
R632 x1.ADJ x2.OUT.t4 53.3636
R633 x2.x2.Z x2.OUT.t0 41.6352
R634 x2.x2.Z x1.ADJ 6.3988
R635 x2.x2.Z x2.OUT.t2 1.35076
R636 EN_N.n2 EN_N.t3 1043.05
R637 EN_N.t3 EN_N.n1 1040.82
R638 EN_N.n1 EN_N.t1 194.654
R639 EN_N.n3 EN_N.t2 7.78263
R640 EN_N.n4 EN_N.t0 6.12265
R641 EN_N.n4 EN_N.n3 2.50721
R642 EN_N.n0 EN_N 1.72738
R643 EN_N.n3 EN_N.n2 1.70148
R644 EN_N.n4 EN_N 1.2505
R645 EN_N.n2 EN_N.n0 0.557375
R646 EN_N.n1 EN_N.n0 0.163
R647 EN_N EN_N.n4 0.063
R648 x1.pg2g x1.pg2g.t1 61.169
R649 x1.pg2g x1.pg2g.t2 22.3222
R650 x1.pg2g x1.pg2g.t0 21.7234
R651 RESULT.n6 RESULT.t4 113.796
R652 RESULT.n4 RESULT.t0 84.6387
R653 RESULT.n1 RESULT.t3 61.3556
R654 RESULT.n3 RESULT.t1 41.6943
R655 RESULT RESULT.t2 41.5734
R656 RESULT.n5 RESULT 3.56033
R657 RESULT.n5 RESULT.n4 3.52161
R658 RESULT.n6 RESULT.n5 2.22055
R659 RESULT.n4 RESULT.n3 1.59772
R660 RESULT.n3 RESULT.n2 0.323684
R661 RESULT.n0 RESULT 0.208833
R662 RESULT.n0 RESULT 0.179071
R663 RESULT.n1 RESULT 0.119281
R664 RESULT RESULT.n7 0.0772045
R665 RESULT.n7 RESULT.n0 0.0734167
R666 RESULT.n2 RESULT 0.0587461
R667 RESULT.n7 RESULT.n6 0.03225
R668 RESULT.n2 RESULT.n1 0.0070445
R669 x1.mirhigh.n0 x1.mirhigh.t1 73.9922
R670 x1.mirhigh x1.mirhigh.t2 62.3033
R671 x1.mirhigh.n0 x1.mirhigh.t0 48.1635
R672 x1.mirhigh x1.mirhigh.n0 1.99219
R673 CALIB.n1 CALIB.t0 234.692
R674 CALIB CALIB.t3 233.88
R675 CALIB.n2 CALIB.t6 229.185
R676 CALIB.n7 CALIB.t2 193.226
R677 CALIB.n0 CALIB.t1 193.153
R678 CALIB.n0 CALIB.t4 174.048
R679 CALIB.n8 CALIB.t5 174.005
R680 CALIB.n12 CALIB.n0 12.9781
R681 CALIB.n1 CALIB 4.63738
R682 CALIB.n3 CALIB.n2 4.5005
R683 CALIB.n0 CALIB 1.89741
R684 CALIB.n11 CALIB.n10 1.46824
R685 CALIB.n7 CALIB 1.188
R686 CALIB.n0 CALIB 1.188
R687 CALIB.n10 CALIB.n9 1.10352
R688 CALIB.n9 CALIB.n6 1.09448
R689 CALIB.n3 CALIB 1.04576
R690 CALIB.n9 CALIB.n8 0.853
R691 CALIB.n6 CALIB.n5 0.559652
R692 CALIB.n12 CALIB.n11 0.203625
R693 CALIB.n5 CALIB.n4 0.188
R694 CALIB.n4 CALIB 0.180647
R695 CALIB.n6 CALIB.n2 0.124054
R696 CALIB.n8 CALIB.n7 0.0820074
R697 CALIB CALIB.n12 0.063
R698 CALIB.n11 CALIB 0.041125
R699 CALIB.n10 CALIB.n1 0.0394785
R700 CALIB.n5 CALIB 0.0194732
R701 CALIB.n4 CALIB.n3 0.00481034
C0 x1.pg2g x1.G2 0.153401f
C1 x1.p2p EN_N 0.150607f
C2 x1.G1 THRESHV 1.40388f
C3 VCC x1.n2n 0.200319f
C4 CALIB INPUT 0.941608f
C5 EN_N RESULT 0.916484f
C6 CALIB x2.x2.GP 1.13808f
C7 x3.OUT EN_N 0.040617f
C8 x3.OUT INPUT 0.624154f
C9 CALIB VCC 4.035002f
C10 VCC x1.p2p 0.888453f
C11 x2.x2.GP RESULT 0.976261f
C12 CALIB x1.G2 0.027326f
C13 x1.G1 EN_N 0.15289f
C14 x3.OUT x1.inhigh 0.692478f
C15 VCC RESULT 1.9672f
C16 x1.mirhigh RESULT 0.15303f
C17 VCC x3.OUT 2.816242f
C18 x3.OUT x1.mirhigh 1.41e-19
C19 x1.G2 RESULT 0.471118f
C20 x3.OUT x1.G2 1.28923f
C21 x1.G1 x1.inhigh 0.896861f
C22 EN_N THRESHV 0.235529f
C23 VCC x1.G1 1.4999f
C24 x1.G1 x1.mirhigh 0.00484f
C25 INPUT THRESHV 0.554769f
C26 x1.G1 x1.G2 0.305193f
C27 x1.pg2g RESULT 1.16101f
C28 x3.OUT x1.pg2g 4.49e-19
C29 x1.inhigh THRESHV 0.729549f
C30 VCC THRESHV 1.677724f
C31 x1.G1 x1.pg2g 0.397601f
C32 THRESHV x1.G2 0.036113f
C33 CALIB RESULT 0.472262f
C34 x1.G1 x1.n2n 0.676922f
C35 CALIB x3.OUT 1.35366f
C36 EN_N x1.inhigh 0.891479f
C37 VCC EN_N 11.366099f
C38 x1.mirhigh EN_N 0.736523f
C39 VCC INPUT 0.298341f
C40 EN_N x1.G2 0.004728f
C41 CALIB x1.G1 0.026807f
C42 x1.G1 x1.p2p 0.02214f
C43 THRESHV x1.n2n 0.001596f
C44 VCC x2.x2.GP 1.35537f
C45 VCC x1.inhigh 2.00666f
C46 x1.mirhigh x1.inhigh 0.01694f
C47 x1.G1 RESULT 0.010549f
C48 x1.G1 x3.OUT 0.410051f
C49 x1.inhigh x1.G2 0.104764f
C50 VCC x1.mirhigh 3.92074f
C51 EN_N x1.pg2g 0.022928f
C52 CALIB THRESHV 2.03319f
C53 VCC x1.G2 0.932067f
C54 x1.mirhigh x1.G2 0.001507f
C55 EN_N x1.n2n 0.001021f
C56 x1.pg2g x1.inhigh 0.00845f
C57 x3.OUT THRESHV 1.39678f
C58 VCC x1.pg2g 3.78855f
C59 x1.mirhigh x1.pg2g 1.02871f
C60 x1.inhigh x1.n2n 5.52e-19
C61 INPUT VSS 1.38167f
C62 CALIB VSS 9.496784f
C63 RESULT VSS 6.95466f
C64 THRESHV VSS 5.571935f
C65 EN_N VSS 8.190082f
C66 VCC VSS 65.513626f
C67 x2.x2.GP VSS 0.927891f
C68 x1.pg2g VSS 4.93169f
C69 x1.G2 VSS 9.06897f
C70 x3.OUT VSS 6.915897f
C71 x1.n2n VSS 0.996702f
C72 x1.G1 VSS 7.98487f
C73 x1.mirhigh VSS 1.527153f
C74 x1.inhigh VSS 2.94796f
C75 x1.p2p VSS 0.150606f
C76 CALIB.t1 VSS 0.016344f
C77 CALIB.t4 VSS 0.050439f
C78 CALIB.t3 VSS 0.0313f
C79 CALIB.n0 VSS 2.08039f
C80 CALIB.t0 VSS 0.027969f
C81 CALIB.n1 VSS 0.175296f
C82 CALIB.t6 VSS 0.027457f
C83 CALIB.n2 VSS 0.208588f
C84 CALIB.n3 VSS 0.007374f
C85 CALIB.n4 VSS 0.010406f
C86 CALIB.n5 VSS 0.087216f
C87 CALIB.n6 VSS 0.155746f
C88 CALIB.t5 VSS 0.050387f
C89 CALIB.t2 VSS 0.016421f
C90 CALIB.n7 VSS 0.240185f
C91 CALIB.n8 VSS 0.23243f
C92 CALIB.n9 VSS 0.705296f
C93 CALIB.n10 VSS 0.049017f
C94 CALIB.n11 VSS 0.067385f
C95 CALIB.n12 VSS 0.933453f
C96 x1.mirhigh.t2 VSS 0.241652f
C97 x1.mirhigh.t1 VSS 0.472059f
C98 x1.mirhigh.t0 VSS 0.294208f
C99 x1.mirhigh.n0 VSS 2.23501f
C100 x1.pg2g.t2 VSS 0.771449f
C101 x1.pg2g.t0 VSS 0.738093f
C102 x1.pg2g.t1 VSS 0.060558f
C103 EN_N.t0 VSS 1.29992f
C104 EN_N.n0 VSS 0.59083f
C105 EN_N.t1 VSS 0.045334f
C106 EN_N.n1 VSS 2.42458f
C107 EN_N.t3 VSS 0.05422f
C108 EN_N.n2 VSS 0.986737f
C109 EN_N.t2 VSS 1.84923f
C110 EN_N.n3 VSS 2.4026f
C111 EN_N.n4 VSS 1.56361f
C112 x2.OUT.t2 VSS 1.20129f
C113 x2.x2.Z VSS 0.787408f
C114 x1.ADJ VSS 0.102848f
C115 x2.OUT.t4 VSS 0.002626f
C116 x2.OUT.t3 VSS 0.003534f
C117 x2.OUT.t1 VSS 0.001163f
C118 x2.OUT.t0 VSS 0.001127f
C119 VCC.n0 VSS 0.954377f
C120 VCC.t15 VSS 0.764334f
C121 VCC.n1 VSS 0.024789f
C122 VCC.n2 VSS 0.024901f
C123 VCC.n4 VSS 0.025358f
C124 VCC.n5 VSS 0.025337f
C125 VCC.n6 VSS 0.175596f
C126 VCC.t8 VSS 0.252681f
C127 VCC.n8 VSS 0.025358f
C128 VCC.n9 VSS 0.175596f
C129 VCC.n10 VSS 0.017774f
C130 VCC.n11 VSS 0.017728f
C131 VCC.n12 VSS 0.787446f
C132 VCC.n13 VSS 0.038595f
C133 VCC.n14 VSS 0.031601f
C134 VCC.n15 VSS 0.540291f
C135 VCC.n16 VSS 0.540291f
C136 VCC.n17 VSS 0.036791f
C137 VCC.n18 VSS 0.052501f
C138 VCC.n19 VSS 0.053587f
C139 VCC.n21 VSS 0.055231f
C140 VCC.n22 VSS 0.055222f
C141 VCC.n23 VSS 0.625537f
C142 VCC.t7 VSS 1.02077f
C143 VCC.n25 VSS 0.055231f
C144 VCC.n26 VSS 0.625537f
C145 VCC.n27 VSS 0.045226f
C146 VCC.n28 VSS 0.045615f
C147 VCC.n29 VSS 0.050618f
C148 VCC.n30 VSS 0.065584f
C149 VCC.n32 VSS 0.065584f
C150 VCC.n33 VSS 0.064789f
C151 VCC.n34 VSS 0.706368f
C152 VCC.t9 VSS 1.08096f
C153 VCC.n36 VSS 0.065584f
C154 VCC.n37 VSS 0.706368f
C155 VCC.n38 VSS 0.045885f
C156 VCC.n39 VSS 0.055163f
C157 VCC.n40 VSS 0.614895f
C158 VCC.n41 VSS 0.033838f
C159 VCC.n42 VSS 0.055231f
C160 VCC.n43 VSS 0.055231f
C161 VCC.t10 VSS 1.02077f
C162 VCC.n44 VSS 0.054079f
C163 VCC.n46 VSS 0.625537f
C164 VCC.n47 VSS 0.055231f
C165 VCC.n49 VSS 0.625537f
C166 VCC.n50 VSS 0.05391f
C167 VCC.n51 VSS 0.037528f
C168 VCC.n52 VSS 1.75862f
C169 VCC.t12 VSS 0.078086f
C170 VCC.n53 VSS 0.968801f
C171 VCC.n54 VSS 0.038276f
C172 VCC.n55 VSS 0.040483f
C173 VCC.n56 VSS 0.040483f
C174 VCC.t11 VSS 0.439376f
C175 VCC.n57 VSS 0.044328f
C176 VCC.n59 VSS 0.266303f
C177 VCC.n60 VSS 0.040483f
C178 VCC.n62 VSS 0.266303f
C179 VCC.n63 VSS 0.0444f
C180 VCC.n64 VSS 0.038158f
C181 VCC.n65 VSS 0.742778f
C182 VCC.n66 VSS 0.960922f
C183 VCC.t14 VSS 0.03114f
C184 VCC.n67 VSS 0.037795f
C185 VCC.n68 VSS 0.067947f
C186 VCC.n69 VSS 0.695711f
C187 VCC.n70 VSS 0.695711f
C188 VCC.n71 VSS 0.062643f
C189 VCC.n72 VSS 0.062753f
C190 VCC.n73 VSS 0.064797f
C191 VCC.t13 VSS 1.18469f
C192 VCC.n76 VSS 0.064797f
C193 VCC.n77 VSS 0.06367f
C194 VCC.n78 VSS 0.035773f
C195 VCC.n79 VSS 0.066668f
C196 VCC.n80 VSS 0.045937f
C197 VCC.n81 VSS 0.065584f
C198 VCC.n83 VSS 0.065584f
C199 VCC.n84 VSS 0.064789f
C200 VCC.n85 VSS 0.706368f
C201 VCC.t0 VSS 1.08096f
C202 VCC.n87 VSS 0.065584f
C203 VCC.n88 VSS 0.706368f
C204 VCC.n89 VSS 0.05035f
C205 VCC.n90 VSS 0.064041f
C206 VCC.t6 VSS 0.015618f
C207 VCC.n91 VSS 0.09394f
C208 VCC.n92 VSS 0.35588f
C209 VCC.n93 VSS 0.084052f
C210 VCC.n94 VSS 0.615732f
C211 VCC.n95 VSS 1.14824f
C212 VCC.n96 VSS 0.06798f
C213 VCC.n97 VSS 0.068606f
C214 VCC.n98 VSS 0.059714f
C215 VCC.t5 VSS 0.902255f
C216 VCC.n101 VSS 0.059714f
C217 VCC.n102 VSS 0.0588f
C218 VCC.n103 VSS 0.032602f
C219 VCC.n104 VSS 0.299596f
C220 x1.inhigh.t2 VSS 0.040812f
C221 x1.inhigh.t1 VSS 0.141031f
C222 x1.inhigh.t0 VSS 0.141031f
C223 THRESHV.t1 VSS 0.021224f
C224 THRESHV.t0 VSS 0.020509f
C225 THRESHV.n0 VSS 0.033562f
C226 THRESHV.n1 VSS 0.51856f
C227 THRESHV.n2 VSS 0.289799f
C228 THRESHV.n3 VSS 0.036223f
C229 THRESHV.t2 VSS 0.432963f
C230 THRESHV.n4 VSS 1.4611f
C231 THRESHV.n5 VSS 0.718266f
C232 x3.OUT.n0 VSS 1.19689f
C233 x3.OUT.t3 VSS 0.014249f
C234 x3.OUT.t4 VSS 0.290549f
C235 x3.OUT.t2 VSS 0.013538f
C236 x3.OUT.t1 VSS 0.014256f
C237 x3.OUT.t0 VSS 0.013797f
C238 x3.x2.GP VSS 1.20755f
C239 x3.SEL_N.t3 VSS 0.023118f
C240 x3.SEL_N.t2 VSS 0.023076f
C241 x3.x3.GN VSS 0.807187f
C242 x3.SEL_N.t0 VSS 0.026392f
C243 x3.SEL_N.t1 VSS 0.01268f
.ends

