MACRO p3_opamp
  CLASS BLOCK ;
  FOREIGN p3_opamp ;
  ORIGIN -18.250 -15.850 ;
  SIZE 24.250 BY 25.450 ;
  PIN VDD
    ANTENNADIFFAREA 23.521200 ;
    PORT
      LAYER met1 ;
        RECT 19.900 39.400 20.900 40.400 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 25.696999 ;
    PORT
      LAYER met1 ;
        RECT 19.350 16.550 20.350 17.550 ;
    END
  END VSS
  PIN PLUS
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met1 ;
        RECT 33.250 21.650 34.250 22.650 ;
    END
  END PLUS
  PIN MINUS
    ANTENNAGATEAREA 1.250000 ;
    PORT
      LAYER met1 ;
        RECT 23.400 21.650 24.400 22.650 ;
    END
  END MINUS
  PIN VOUT
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met1 ;
        RECT 39.850 36.200 40.850 37.200 ;
    END
  END VOUT
  OBS
      LAYER pwell ;
        RECT 20.000 29.400 22.010 38.020 ;
        RECT 19.450 17.750 22.550 28.580 ;
      LAYER nwell ;
        RECT 24.050 23.800 27.240 39.210 ;
        RECT 30.400 23.800 33.590 39.210 ;
      LAYER pwell ;
        RECT 24.200 20.950 33.400 23.410 ;
      LAYER nwell ;
        RECT 35.000 22.000 38.190 39.470 ;
      LAYER pwell ;
        RECT 31.000 20.900 31.550 20.950 ;
        RECT 23.500 17.800 34.330 20.900 ;
        RECT 39.000 17.800 42.100 35.500 ;
      LAYER li1 ;
        RECT 35.180 39.120 38.010 39.290 ;
        RECT 24.230 38.860 27.060 39.030 ;
        RECT 24.230 38.500 24.400 38.860 ;
        RECT 20.180 37.670 21.830 37.840 ;
        RECT 20.180 37.350 20.350 37.670 ;
        RECT 20.100 30.200 20.350 37.350 ;
        RECT 20.830 35.030 21.180 37.190 ;
        RECT 20.830 30.230 21.180 32.390 ;
        RECT 20.180 29.750 20.350 30.200 ;
        RECT 21.660 29.750 21.830 37.670 ;
        RECT 20.180 29.580 21.830 29.750 ;
        RECT 19.630 28.300 22.370 28.400 ;
        RECT 19.550 28.230 22.370 28.300 ;
        RECT 19.550 18.950 19.800 28.230 ;
        RECT 20.480 27.660 21.520 27.830 ;
        RECT 20.140 25.600 20.310 27.600 ;
        RECT 21.690 25.600 21.860 27.600 ;
        RECT 20.480 25.370 21.520 25.540 ;
        RECT 20.140 23.310 20.310 25.310 ;
        RECT 21.690 23.310 21.860 25.310 ;
        RECT 20.480 23.080 21.520 23.250 ;
        RECT 20.140 21.020 20.310 23.020 ;
        RECT 21.690 21.020 21.860 23.020 ;
        RECT 20.480 20.790 21.520 20.960 ;
        RECT 19.630 18.100 19.800 18.950 ;
        RECT 20.140 18.730 20.310 20.730 ;
        RECT 21.690 18.730 21.860 20.730 ;
        RECT 20.480 18.500 21.520 18.670 ;
        RECT 20.050 18.100 21.950 18.150 ;
        RECT 22.200 18.100 22.370 28.230 ;
        RECT 24.100 26.600 24.400 38.500 ;
        RECT 25.125 38.290 26.165 38.460 ;
        RECT 24.740 36.230 24.910 38.230 ;
        RECT 26.380 36.230 26.550 38.230 ;
        RECT 25.125 36.000 26.165 36.170 ;
        RECT 24.740 33.940 24.910 35.940 ;
        RECT 26.380 33.940 26.550 35.940 ;
        RECT 25.125 33.710 26.165 33.880 ;
        RECT 24.740 31.650 24.910 33.650 ;
        RECT 26.380 31.650 26.550 33.650 ;
        RECT 25.125 31.420 26.165 31.590 ;
        RECT 24.740 29.360 24.910 31.360 ;
        RECT 26.380 29.360 26.550 31.360 ;
        RECT 25.125 29.130 26.165 29.300 ;
        RECT 24.740 27.070 24.910 29.070 ;
        RECT 26.380 27.070 26.550 29.070 ;
        RECT 25.125 26.840 26.165 27.010 ;
        RECT 24.230 24.150 24.400 26.600 ;
        RECT 24.740 24.780 24.910 26.780 ;
        RECT 26.380 24.780 26.550 26.780 ;
        RECT 25.125 24.550 26.165 24.720 ;
        RECT 26.890 24.150 27.060 38.860 ;
        RECT 24.230 23.980 27.060 24.150 ;
        RECT 30.580 38.860 33.410 39.030 ;
        RECT 30.580 24.150 30.750 38.860 ;
        RECT 33.240 38.500 33.410 38.860 ;
        RECT 35.180 38.750 35.350 39.120 ;
        RECT 31.475 38.290 32.515 38.460 ;
        RECT 31.090 36.230 31.260 38.230 ;
        RECT 32.730 36.230 32.900 38.230 ;
        RECT 31.475 36.000 32.515 36.170 ;
        RECT 31.090 33.940 31.260 35.940 ;
        RECT 32.730 33.940 32.900 35.940 ;
        RECT 31.475 33.710 32.515 33.880 ;
        RECT 31.090 31.650 31.260 33.650 ;
        RECT 32.730 31.650 32.900 33.650 ;
        RECT 31.475 31.420 32.515 31.590 ;
        RECT 31.090 29.360 31.260 31.360 ;
        RECT 32.730 29.360 32.900 31.360 ;
        RECT 31.475 29.130 32.515 29.300 ;
        RECT 31.090 27.070 31.260 29.070 ;
        RECT 32.730 27.070 32.900 29.070 ;
        RECT 31.475 26.840 32.515 27.010 ;
        RECT 31.090 24.780 31.260 26.780 ;
        RECT 32.730 24.780 32.900 26.780 ;
        RECT 33.240 26.600 33.550 38.500 ;
        RECT 31.475 24.550 32.515 24.720 ;
        RECT 33.240 24.150 33.410 26.600 ;
        RECT 30.580 23.980 33.410 24.150 ;
        RECT 24.380 23.060 28.620 23.230 ;
        RECT 24.380 21.300 24.550 23.060 ;
        RECT 25.230 22.490 27.770 22.660 ;
        RECT 24.890 21.930 25.060 22.430 ;
        RECT 27.940 21.930 28.110 22.430 ;
        RECT 25.230 21.700 27.770 21.870 ;
        RECT 28.450 21.300 28.620 23.060 ;
        RECT 24.380 21.130 28.620 21.300 ;
        RECT 28.980 23.060 33.220 23.230 ;
        RECT 35.150 23.200 35.350 38.750 ;
        RECT 36.075 38.550 37.115 38.720 ;
        RECT 35.690 37.990 35.860 38.490 ;
        RECT 37.330 37.990 37.500 38.490 ;
        RECT 36.075 37.760 37.115 37.930 ;
        RECT 35.690 37.200 35.860 37.700 ;
        RECT 37.330 37.200 37.500 37.700 ;
        RECT 36.075 36.970 37.115 37.140 ;
        RECT 35.690 36.410 35.860 36.910 ;
        RECT 37.330 36.410 37.500 36.910 ;
        RECT 36.075 36.180 37.115 36.350 ;
        RECT 35.690 35.620 35.860 36.120 ;
        RECT 37.330 35.620 37.500 36.120 ;
        RECT 36.075 35.390 37.115 35.560 ;
        RECT 35.690 34.830 35.860 35.330 ;
        RECT 37.330 34.830 37.500 35.330 ;
        RECT 36.075 34.600 37.115 34.770 ;
        RECT 35.690 34.040 35.860 34.540 ;
        RECT 37.330 34.040 37.500 34.540 ;
        RECT 36.075 33.810 37.115 33.980 ;
        RECT 35.690 33.250 35.860 33.750 ;
        RECT 37.330 33.250 37.500 33.750 ;
        RECT 36.075 33.020 37.115 33.190 ;
        RECT 35.690 32.460 35.860 32.960 ;
        RECT 37.330 32.460 37.500 32.960 ;
        RECT 36.075 32.230 37.115 32.400 ;
        RECT 35.690 31.670 35.860 32.170 ;
        RECT 37.330 31.670 37.500 32.170 ;
        RECT 36.075 31.440 37.115 31.610 ;
        RECT 35.690 30.880 35.860 31.380 ;
        RECT 37.330 30.880 37.500 31.380 ;
        RECT 36.075 30.650 37.115 30.820 ;
        RECT 35.690 30.090 35.860 30.590 ;
        RECT 37.330 30.090 37.500 30.590 ;
        RECT 36.075 29.860 37.115 30.030 ;
        RECT 35.690 29.300 35.860 29.800 ;
        RECT 37.330 29.300 37.500 29.800 ;
        RECT 36.075 29.070 37.115 29.240 ;
        RECT 35.690 28.510 35.860 29.010 ;
        RECT 37.330 28.510 37.500 29.010 ;
        RECT 36.075 28.280 37.115 28.450 ;
        RECT 35.690 27.720 35.860 28.220 ;
        RECT 37.330 27.720 37.500 28.220 ;
        RECT 36.075 27.490 37.115 27.660 ;
        RECT 35.690 26.930 35.860 27.430 ;
        RECT 37.330 26.930 37.500 27.430 ;
        RECT 36.075 26.700 37.115 26.870 ;
        RECT 35.690 26.140 35.860 26.640 ;
        RECT 37.330 26.140 37.500 26.640 ;
        RECT 36.075 25.910 37.115 26.080 ;
        RECT 35.690 25.350 35.860 25.850 ;
        RECT 37.330 25.350 37.500 25.850 ;
        RECT 36.075 25.120 37.115 25.290 ;
        RECT 35.690 24.560 35.860 25.060 ;
        RECT 37.330 24.560 37.500 25.060 ;
        RECT 36.075 24.330 37.115 24.500 ;
        RECT 35.690 23.770 35.860 24.270 ;
        RECT 37.330 23.770 37.500 24.270 ;
        RECT 36.075 23.540 37.115 23.710 ;
        RECT 28.980 21.300 29.150 23.060 ;
        RECT 29.830 22.490 32.370 22.660 ;
        RECT 29.490 21.930 29.660 22.430 ;
        RECT 32.540 21.930 32.710 22.430 ;
        RECT 29.830 21.700 32.370 21.870 ;
        RECT 33.050 21.300 33.220 23.060 ;
        RECT 35.180 22.350 35.350 23.200 ;
        RECT 35.690 22.980 35.860 23.480 ;
        RECT 37.330 22.980 37.500 23.480 ;
        RECT 36.075 22.750 37.115 22.920 ;
        RECT 37.840 22.350 38.010 39.120 ;
        RECT 35.180 22.180 38.010 22.350 ;
        RECT 39.180 35.150 41.920 35.320 ;
        RECT 28.980 21.130 33.350 21.300 ;
        RECT 24.400 21.100 25.200 21.130 ;
        RECT 32.550 21.100 33.350 21.130 ;
        RECT 19.630 17.930 22.370 18.100 ;
        RECT 23.680 20.550 34.150 20.720 ;
        RECT 23.680 18.150 23.850 20.550 ;
        RECT 24.480 20.040 26.480 20.210 ;
        RECT 26.770 20.040 28.770 20.210 ;
        RECT 29.060 20.040 31.060 20.210 ;
        RECT 31.350 20.040 33.350 20.210 ;
        RECT 33.980 20.050 34.150 20.550 ;
        RECT 24.250 18.830 24.420 19.870 ;
        RECT 26.540 18.830 26.710 19.870 ;
        RECT 28.830 18.830 29.000 19.870 ;
        RECT 31.120 18.830 31.290 19.870 ;
        RECT 33.410 18.830 33.580 19.870 ;
        RECT 24.480 18.490 26.480 18.660 ;
        RECT 26.770 18.490 28.770 18.660 ;
        RECT 29.060 18.490 31.060 18.660 ;
        RECT 31.350 18.490 33.350 18.660 ;
        RECT 33.950 18.450 34.200 20.050 ;
        RECT 39.180 19.600 39.350 35.150 ;
        RECT 40.030 34.580 41.070 34.750 ;
        RECT 39.690 32.520 39.860 34.520 ;
        RECT 41.240 32.520 41.410 34.520 ;
        RECT 40.030 32.290 41.070 32.460 ;
        RECT 39.690 30.230 39.860 32.230 ;
        RECT 41.240 30.230 41.410 32.230 ;
        RECT 40.030 30.000 41.070 30.170 ;
        RECT 39.690 27.940 39.860 29.940 ;
        RECT 41.240 27.940 41.410 29.940 ;
        RECT 40.030 27.710 41.070 27.880 ;
        RECT 39.690 25.650 39.860 27.650 ;
        RECT 41.240 25.650 41.410 27.650 ;
        RECT 40.030 25.420 41.070 25.590 ;
        RECT 39.690 23.360 39.860 25.360 ;
        RECT 41.240 23.360 41.410 25.360 ;
        RECT 40.030 23.130 41.070 23.300 ;
        RECT 39.690 21.070 39.860 23.070 ;
        RECT 41.240 21.070 41.410 23.070 ;
        RECT 40.030 20.840 41.070 21.010 ;
        RECT 39.100 18.450 39.350 19.600 ;
        RECT 39.690 18.780 39.860 20.780 ;
        RECT 41.240 18.780 41.410 20.780 ;
        RECT 41.750 19.600 41.920 35.150 ;
        RECT 40.030 18.550 41.070 18.720 ;
        RECT 33.980 18.150 34.150 18.450 ;
        RECT 23.680 17.980 34.150 18.150 ;
        RECT 39.180 18.150 39.350 18.450 ;
        RECT 41.750 18.450 42.000 19.600 ;
        RECT 41.750 18.150 41.920 18.450 ;
        RECT 39.180 17.980 41.920 18.150 ;
        RECT 20.050 17.850 21.950 17.930 ;
        RECT 24.150 17.900 33.700 17.980 ;
        RECT 39.450 17.950 41.650 17.980 ;
      LAYER mcon ;
        RECT 20.100 30.200 20.350 37.350 ;
        RECT 20.910 35.115 21.100 37.100 ;
        RECT 20.910 30.320 21.100 32.305 ;
        RECT 19.550 18.950 19.800 28.300 ;
        RECT 20.560 27.660 21.440 27.830 ;
        RECT 20.140 25.680 20.310 27.520 ;
        RECT 21.690 25.680 21.860 27.520 ;
        RECT 20.560 25.370 21.440 25.540 ;
        RECT 20.140 23.390 20.310 25.230 ;
        RECT 21.690 23.390 21.860 25.230 ;
        RECT 20.560 23.080 21.440 23.250 ;
        RECT 20.140 21.100 20.310 22.940 ;
        RECT 21.690 21.100 21.860 22.940 ;
        RECT 20.560 20.790 21.440 20.960 ;
        RECT 20.140 18.810 20.310 20.650 ;
        RECT 21.690 18.810 21.860 20.650 ;
        RECT 20.560 18.500 21.440 18.670 ;
        RECT 24.100 26.600 24.400 38.500 ;
        RECT 25.205 38.290 26.085 38.460 ;
        RECT 24.740 36.310 24.910 38.150 ;
        RECT 26.380 36.310 26.550 38.150 ;
        RECT 25.205 36.000 26.085 36.170 ;
        RECT 24.740 34.020 24.910 35.860 ;
        RECT 26.380 34.020 26.550 35.860 ;
        RECT 25.205 33.710 26.085 33.880 ;
        RECT 24.740 31.730 24.910 33.570 ;
        RECT 26.380 31.730 26.550 33.570 ;
        RECT 25.205 31.420 26.085 31.590 ;
        RECT 24.740 29.440 24.910 31.280 ;
        RECT 26.380 29.440 26.550 31.280 ;
        RECT 25.205 29.130 26.085 29.300 ;
        RECT 24.740 27.150 24.910 28.990 ;
        RECT 26.380 27.150 26.550 28.990 ;
        RECT 25.205 26.840 26.085 27.010 ;
        RECT 24.740 24.860 24.910 26.700 ;
        RECT 26.380 24.860 26.550 26.700 ;
        RECT 25.205 24.550 26.085 24.720 ;
        RECT 31.555 38.290 32.435 38.460 ;
        RECT 31.090 36.310 31.260 38.150 ;
        RECT 32.730 36.310 32.900 38.150 ;
        RECT 31.555 36.000 32.435 36.170 ;
        RECT 31.090 34.020 31.260 35.860 ;
        RECT 32.730 34.020 32.900 35.860 ;
        RECT 31.555 33.710 32.435 33.880 ;
        RECT 31.090 31.730 31.260 33.570 ;
        RECT 32.730 31.730 32.900 33.570 ;
        RECT 31.555 31.420 32.435 31.590 ;
        RECT 31.090 29.440 31.260 31.280 ;
        RECT 32.730 29.440 32.900 31.280 ;
        RECT 31.555 29.130 32.435 29.300 ;
        RECT 31.090 27.150 31.260 28.990 ;
        RECT 32.730 27.150 32.900 28.990 ;
        RECT 31.555 26.840 32.435 27.010 ;
        RECT 31.090 24.860 31.260 26.700 ;
        RECT 32.730 24.860 32.900 26.700 ;
        RECT 33.250 26.600 33.550 38.500 ;
        RECT 31.555 24.550 32.435 24.720 ;
        RECT 25.310 22.490 27.690 22.660 ;
        RECT 24.890 22.010 25.060 22.350 ;
        RECT 27.940 22.010 28.110 22.350 ;
        RECT 25.310 21.700 27.690 21.870 ;
        RECT 35.150 23.200 35.350 38.750 ;
        RECT 36.155 38.550 37.035 38.720 ;
        RECT 35.690 38.070 35.860 38.410 ;
        RECT 37.330 38.070 37.500 38.410 ;
        RECT 36.155 37.760 37.035 37.930 ;
        RECT 35.690 37.280 35.860 37.620 ;
        RECT 37.330 37.280 37.500 37.620 ;
        RECT 36.155 36.970 37.035 37.140 ;
        RECT 35.690 36.490 35.860 36.830 ;
        RECT 37.330 36.490 37.500 36.830 ;
        RECT 36.155 36.180 37.035 36.350 ;
        RECT 35.690 35.700 35.860 36.040 ;
        RECT 37.330 35.700 37.500 36.040 ;
        RECT 36.155 35.390 37.035 35.560 ;
        RECT 35.690 34.910 35.860 35.250 ;
        RECT 37.330 34.910 37.500 35.250 ;
        RECT 36.155 34.600 37.035 34.770 ;
        RECT 35.690 34.120 35.860 34.460 ;
        RECT 37.330 34.120 37.500 34.460 ;
        RECT 36.155 33.810 37.035 33.980 ;
        RECT 35.690 33.330 35.860 33.670 ;
        RECT 37.330 33.330 37.500 33.670 ;
        RECT 36.155 33.020 37.035 33.190 ;
        RECT 35.690 32.540 35.860 32.880 ;
        RECT 37.330 32.540 37.500 32.880 ;
        RECT 36.155 32.230 37.035 32.400 ;
        RECT 35.690 31.750 35.860 32.090 ;
        RECT 37.330 31.750 37.500 32.090 ;
        RECT 36.155 31.440 37.035 31.610 ;
        RECT 35.690 30.960 35.860 31.300 ;
        RECT 37.330 30.960 37.500 31.300 ;
        RECT 36.155 30.650 37.035 30.820 ;
        RECT 35.690 30.170 35.860 30.510 ;
        RECT 37.330 30.170 37.500 30.510 ;
        RECT 36.155 29.860 37.035 30.030 ;
        RECT 35.690 29.380 35.860 29.720 ;
        RECT 37.330 29.380 37.500 29.720 ;
        RECT 36.155 29.070 37.035 29.240 ;
        RECT 35.690 28.590 35.860 28.930 ;
        RECT 37.330 28.590 37.500 28.930 ;
        RECT 36.155 28.280 37.035 28.450 ;
        RECT 35.690 27.800 35.860 28.140 ;
        RECT 37.330 27.800 37.500 28.140 ;
        RECT 36.155 27.490 37.035 27.660 ;
        RECT 35.690 27.010 35.860 27.350 ;
        RECT 37.330 27.010 37.500 27.350 ;
        RECT 36.155 26.700 37.035 26.870 ;
        RECT 35.690 26.220 35.860 26.560 ;
        RECT 37.330 26.220 37.500 26.560 ;
        RECT 36.155 25.910 37.035 26.080 ;
        RECT 35.690 25.430 35.860 25.770 ;
        RECT 37.330 25.430 37.500 25.770 ;
        RECT 36.155 25.120 37.035 25.290 ;
        RECT 35.690 24.640 35.860 24.980 ;
        RECT 37.330 24.640 37.500 24.980 ;
        RECT 36.155 24.330 37.035 24.500 ;
        RECT 35.690 23.850 35.860 24.190 ;
        RECT 37.330 23.850 37.500 24.190 ;
        RECT 36.155 23.540 37.035 23.710 ;
        RECT 29.910 22.490 32.290 22.660 ;
        RECT 29.490 22.010 29.660 22.350 ;
        RECT 32.540 22.010 32.710 22.350 ;
        RECT 29.910 21.700 32.290 21.870 ;
        RECT 35.690 23.060 35.860 23.400 ;
        RECT 37.330 23.060 37.500 23.400 ;
        RECT 36.155 22.750 37.035 22.920 ;
        RECT 24.560 20.040 26.400 20.210 ;
        RECT 26.850 20.040 28.690 20.210 ;
        RECT 29.140 20.040 30.980 20.210 ;
        RECT 31.430 20.040 33.270 20.210 ;
        RECT 24.250 18.910 24.420 19.790 ;
        RECT 26.540 18.910 26.710 19.790 ;
        RECT 28.830 18.910 29.000 19.790 ;
        RECT 31.120 18.910 31.290 19.790 ;
        RECT 33.410 18.910 33.580 19.790 ;
        RECT 24.560 18.490 26.400 18.660 ;
        RECT 26.850 18.490 28.690 18.660 ;
        RECT 29.140 18.490 30.980 18.660 ;
        RECT 31.430 18.490 33.270 18.660 ;
        RECT 40.110 34.580 40.990 34.750 ;
        RECT 39.690 32.600 39.860 34.440 ;
        RECT 41.240 32.600 41.410 34.440 ;
        RECT 40.110 32.290 40.990 32.460 ;
        RECT 39.690 30.310 39.860 32.150 ;
        RECT 41.240 30.310 41.410 32.150 ;
        RECT 40.110 30.000 40.990 30.170 ;
        RECT 39.690 28.020 39.860 29.860 ;
        RECT 41.240 28.020 41.410 29.860 ;
        RECT 40.110 27.710 40.990 27.880 ;
        RECT 39.690 25.730 39.860 27.570 ;
        RECT 41.240 25.730 41.410 27.570 ;
        RECT 40.110 25.420 40.990 25.590 ;
        RECT 39.690 23.440 39.860 25.280 ;
        RECT 41.240 23.440 41.410 25.280 ;
        RECT 40.110 23.130 40.990 23.300 ;
        RECT 39.690 21.150 39.860 22.990 ;
        RECT 41.240 21.150 41.410 22.990 ;
        RECT 40.110 20.840 40.990 21.010 ;
        RECT 39.690 18.860 39.860 20.700 ;
        RECT 41.240 18.860 41.410 20.700 ;
        RECT 40.110 18.550 40.990 18.720 ;
      LAYER met1 ;
        RECT 18.250 40.400 42.500 41.300 ;
        RECT 18.250 39.400 19.900 40.400 ;
        RECT 20.900 39.400 42.500 40.400 ;
        RECT 18.250 38.950 42.500 39.400 ;
        RECT 18.250 30.050 20.450 37.800 ;
        RECT 20.600 35.050 21.550 38.950 ;
        RECT 20.880 32.350 21.130 32.365 ;
        RECT 18.250 18.200 19.900 30.050 ;
        RECT 20.750 29.850 22.600 32.350 ;
        RECT 20.500 27.600 21.500 27.950 ;
        RECT 20.110 27.150 20.340 27.580 ;
        RECT 21.650 27.150 22.600 29.850 ;
        RECT 20.100 26.000 22.600 27.150 ;
        RECT 22.750 26.450 24.500 38.950 ;
        RECT 25.100 38.250 30.450 38.600 ;
        RECT 31.450 38.250 32.550 38.550 ;
        RECT 24.710 37.850 24.940 38.210 ;
        RECT 26.300 38.200 30.450 38.250 ;
        RECT 26.300 37.850 30.800 38.200 ;
        RECT 31.060 37.850 31.290 38.210 ;
        RECT 32.700 37.850 32.930 38.210 ;
        RECT 24.700 37.050 32.930 37.850 ;
        RECT 24.700 36.650 28.300 37.050 ;
        RECT 24.710 36.250 24.940 36.650 ;
        RECT 26.300 36.600 28.300 36.650 ;
        RECT 26.350 36.250 28.300 36.600 ;
        RECT 25.150 36.200 26.150 36.250 ;
        RECT 25.145 35.970 26.150 36.200 ;
        RECT 25.150 35.950 26.150 35.970 ;
        RECT 26.400 35.920 28.300 36.250 ;
        RECT 24.710 35.500 24.940 35.920 ;
        RECT 26.350 35.500 28.300 35.920 ;
        RECT 24.700 34.250 28.300 35.500 ;
        RECT 24.710 33.960 24.940 34.250 ;
        RECT 26.300 33.950 28.300 34.250 ;
        RECT 25.100 33.650 28.300 33.950 ;
        RECT 24.710 33.350 24.940 33.630 ;
        RECT 26.300 33.350 28.300 33.650 ;
        RECT 24.700 32.150 28.300 33.350 ;
        RECT 24.710 31.670 24.940 32.150 ;
        RECT 25.150 31.620 26.150 31.650 ;
        RECT 25.145 31.390 26.150 31.620 ;
        RECT 25.150 31.350 26.150 31.390 ;
        RECT 24.710 31.050 24.940 31.340 ;
        RECT 26.300 31.050 28.300 32.150 ;
        RECT 24.700 29.850 28.300 31.050 ;
        RECT 24.710 29.380 24.940 29.850 ;
        RECT 26.300 29.350 28.300 29.850 ;
        RECT 25.100 29.100 28.300 29.350 ;
        RECT 24.710 28.650 24.940 29.050 ;
        RECT 26.300 28.650 28.300 29.100 ;
        RECT 24.700 27.450 28.300 28.650 ;
        RECT 24.710 27.090 24.940 27.450 ;
        RECT 25.150 27.040 26.150 27.100 ;
        RECT 25.145 26.810 26.150 27.040 ;
        RECT 25.150 26.800 26.150 26.810 ;
        RECT 24.710 26.400 24.940 26.760 ;
        RECT 26.300 26.400 28.300 27.450 ;
        RECT 20.110 25.620 20.340 26.000 ;
        RECT 21.650 25.600 22.600 26.000 ;
        RECT 20.500 25.300 22.600 25.600 ;
        RECT 20.110 24.900 20.340 25.290 ;
        RECT 21.650 24.900 22.600 25.300 ;
        RECT 24.700 25.200 28.300 26.400 ;
        RECT 20.100 23.750 22.600 24.900 ;
        RECT 24.710 24.800 24.940 25.200 ;
        RECT 26.300 24.750 28.300 25.200 ;
        RECT 25.100 24.550 28.300 24.750 ;
        RECT 29.300 36.650 32.930 37.050 ;
        RECT 29.300 35.450 30.800 36.650 ;
        RECT 31.060 36.250 31.290 36.650 ;
        RECT 32.700 36.250 32.930 36.650 ;
        RECT 31.500 36.200 32.550 36.250 ;
        RECT 31.495 35.970 32.550 36.200 ;
        RECT 31.500 35.950 32.550 35.970 ;
        RECT 31.060 35.450 31.290 35.920 ;
        RECT 32.700 35.450 32.930 35.920 ;
        RECT 29.300 34.250 32.930 35.450 ;
        RECT 29.300 33.350 30.800 34.250 ;
        RECT 31.060 33.960 31.290 34.250 ;
        RECT 32.700 33.960 32.930 34.250 ;
        RECT 31.450 33.650 32.550 33.950 ;
        RECT 31.060 33.350 31.290 33.630 ;
        RECT 32.700 33.350 32.930 33.630 ;
        RECT 29.300 32.150 32.930 33.350 ;
        RECT 29.300 31.050 30.800 32.150 ;
        RECT 31.060 31.670 31.290 32.150 ;
        RECT 32.700 31.670 32.930 32.150 ;
        RECT 31.500 31.620 32.550 31.650 ;
        RECT 31.495 31.390 32.550 31.620 ;
        RECT 31.500 31.350 32.550 31.390 ;
        RECT 31.060 31.050 31.290 31.340 ;
        RECT 32.700 31.050 32.930 31.340 ;
        RECT 29.300 29.850 32.930 31.050 ;
        RECT 29.300 28.650 30.800 29.850 ;
        RECT 31.060 29.380 31.290 29.850 ;
        RECT 32.700 29.380 32.930 29.850 ;
        RECT 31.450 29.050 32.550 29.350 ;
        RECT 31.060 28.650 31.290 29.050 ;
        RECT 32.700 28.650 32.930 29.050 ;
        RECT 29.300 27.450 32.930 28.650 ;
        RECT 29.300 26.400 30.800 27.450 ;
        RECT 31.060 27.090 31.290 27.450 ;
        RECT 31.500 27.040 32.550 27.100 ;
        RECT 32.700 27.090 32.930 27.450 ;
        RECT 31.495 26.810 32.550 27.040 ;
        RECT 31.500 26.800 32.550 26.810 ;
        RECT 31.060 26.400 31.290 26.760 ;
        RECT 32.700 26.400 32.930 26.760 ;
        RECT 33.100 26.450 35.400 38.950 ;
        RECT 36.050 38.500 37.100 38.800 ;
        RECT 29.300 25.200 32.930 26.400 ;
        RECT 29.300 24.550 30.800 25.200 ;
        RECT 31.060 24.800 31.290 25.200 ;
        RECT 32.700 24.800 32.930 25.200 ;
        RECT 31.775 24.750 32.325 24.780 ;
        RECT 25.100 24.500 30.800 24.550 ;
        RECT 20.110 23.330 20.340 23.750 ;
        RECT 20.500 23.000 21.500 23.350 ;
        RECT 20.110 22.600 20.340 23.000 ;
        RECT 21.650 22.600 22.600 23.750 ;
        RECT 26.300 23.600 30.800 24.500 ;
        RECT 31.450 24.450 32.550 24.750 ;
        RECT 31.550 24.200 32.500 24.450 ;
        RECT 31.775 24.170 32.325 24.200 ;
        RECT 26.300 22.800 28.650 23.600 ;
        RECT 31.500 23.100 32.500 23.500 ;
        RECT 25.400 22.690 28.650 22.800 ;
        RECT 29.950 22.850 32.500 23.100 ;
        RECT 29.950 22.690 32.350 22.850 ;
        RECT 33.550 22.800 35.400 26.450 ;
        RECT 35.550 25.700 35.900 38.500 ;
        RECT 37.300 38.010 37.530 38.470 ;
        RECT 36.100 37.960 37.150 38.000 ;
        RECT 36.095 37.730 37.150 37.960 ;
        RECT 36.100 37.700 37.150 37.730 ;
        RECT 37.300 37.220 37.530 37.680 ;
        RECT 37.900 37.200 42.500 38.050 ;
        RECT 36.050 36.900 37.100 37.200 ;
        RECT 37.300 36.430 37.530 36.890 ;
        RECT 36.100 36.380 37.150 36.400 ;
        RECT 36.095 36.150 37.150 36.380 ;
        RECT 36.100 36.100 37.150 36.150 ;
        RECT 37.900 36.200 39.850 37.200 ;
        RECT 40.850 36.200 42.500 37.200 ;
        RECT 36.050 35.350 37.100 35.650 ;
        RECT 37.300 35.640 37.530 36.100 ;
        RECT 37.300 34.850 37.530 35.310 ;
        RECT 37.900 34.850 42.500 36.200 ;
        RECT 36.100 34.800 37.150 34.850 ;
        RECT 36.095 34.570 37.150 34.800 ;
        RECT 36.100 34.550 37.150 34.570 ;
        RECT 37.900 34.800 41.250 34.850 ;
        RECT 37.300 34.060 37.530 34.520 ;
        RECT 36.050 33.750 37.100 34.050 ;
        RECT 37.300 33.270 37.530 33.730 ;
        RECT 36.100 33.220 37.150 33.250 ;
        RECT 36.095 32.990 37.150 33.220 ;
        RECT 36.100 32.950 37.150 32.990 ;
        RECT 37.300 32.480 37.530 32.940 ;
        RECT 36.050 32.150 37.100 32.450 ;
        RECT 37.300 31.690 37.530 32.150 ;
        RECT 36.100 31.640 37.150 31.650 ;
        RECT 36.095 31.410 37.150 31.640 ;
        RECT 36.100 31.350 37.150 31.410 ;
        RECT 37.300 30.900 37.530 31.360 ;
        RECT 36.050 30.600 37.100 30.900 ;
        RECT 37.300 30.110 37.530 30.570 ;
        RECT 36.100 30.060 37.150 30.100 ;
        RECT 36.095 29.830 37.150 30.060 ;
        RECT 36.100 29.800 37.150 29.830 ;
        RECT 37.300 29.320 37.530 29.780 ;
        RECT 36.050 29.000 37.100 29.300 ;
        RECT 36.100 28.480 37.150 28.550 ;
        RECT 37.300 28.530 37.530 28.990 ;
        RECT 36.095 28.250 37.150 28.480 ;
        RECT 36.050 27.450 37.100 27.750 ;
        RECT 37.300 27.740 37.530 28.200 ;
        RECT 37.300 26.950 37.530 27.410 ;
        RECT 36.100 26.900 37.150 26.950 ;
        RECT 36.095 26.670 37.150 26.900 ;
        RECT 36.100 26.650 37.150 26.670 ;
        RECT 37.300 26.160 37.530 26.620 ;
        RECT 36.050 25.850 37.100 26.150 ;
        RECT 35.550 24.800 35.950 25.700 ;
        RECT 37.300 25.370 37.530 25.830 ;
        RECT 36.100 25.320 37.150 25.350 ;
        RECT 36.095 25.090 37.150 25.320 ;
        RECT 36.100 25.050 37.150 25.090 ;
        RECT 35.550 22.950 35.900 24.800 ;
        RECT 37.300 24.580 37.530 25.040 ;
        RECT 36.050 24.250 37.100 24.550 ;
        RECT 36.100 23.740 37.150 23.800 ;
        RECT 37.300 23.790 37.530 24.250 ;
        RECT 36.095 23.510 37.150 23.740 ;
        RECT 36.100 23.500 37.150 23.510 ;
        RECT 37.300 23.000 37.530 23.460 ;
        RECT 36.050 22.700 37.100 23.000 ;
        RECT 20.100 21.450 22.600 22.600 ;
        RECT 25.250 22.550 28.650 22.690 ;
        RECT 25.250 22.460 27.750 22.550 ;
        RECT 29.850 22.460 32.350 22.690 ;
        RECT 25.400 22.450 27.700 22.460 ;
        RECT 24.860 22.350 25.090 22.410 ;
        RECT 27.910 22.350 28.140 22.410 ;
        RECT 29.460 22.350 29.690 22.410 ;
        RECT 32.510 22.350 32.740 22.410 ;
        RECT 24.750 22.260 25.150 22.350 ;
        RECT 27.850 22.260 28.250 22.350 ;
        RECT 24.400 22.045 28.250 22.260 ;
        RECT 24.750 22.000 25.150 22.045 ;
        RECT 27.850 22.000 28.250 22.045 ;
        RECT 29.350 22.275 29.750 22.350 ;
        RECT 32.450 22.275 32.850 22.350 ;
        RECT 29.350 22.050 33.250 22.275 ;
        RECT 29.350 22.000 29.750 22.050 ;
        RECT 32.450 22.030 33.250 22.050 ;
        RECT 32.450 22.000 32.850 22.030 ;
        RECT 37.900 22.000 39.200 34.800 ;
        RECT 40.000 34.650 41.050 34.800 ;
        RECT 40.050 34.550 41.050 34.650 ;
        RECT 39.660 34.150 39.890 34.500 ;
        RECT 39.550 33.950 39.900 34.150 ;
        RECT 41.210 33.950 41.440 34.500 ;
        RECT 39.550 33.000 41.440 33.950 ;
        RECT 39.550 31.700 39.900 33.000 ;
        RECT 40.050 32.250 41.050 32.550 ;
        RECT 41.210 32.540 41.440 33.000 ;
        RECT 41.210 31.700 41.440 32.210 ;
        RECT 39.550 30.750 41.440 31.700 ;
        RECT 39.550 29.350 39.900 30.750 ;
        RECT 41.210 30.250 41.440 30.750 ;
        RECT 40.050 29.950 41.050 30.250 ;
        RECT 41.210 29.350 41.440 29.920 ;
        RECT 39.550 28.400 41.440 29.350 ;
        RECT 39.550 27.200 39.900 28.400 ;
        RECT 41.210 27.960 41.440 28.400 ;
        RECT 40.050 27.650 41.050 27.950 ;
        RECT 41.210 27.200 41.440 27.630 ;
        RECT 39.550 26.250 41.440 27.200 ;
        RECT 39.550 24.900 39.900 26.250 ;
        RECT 40.050 25.350 41.050 25.700 ;
        RECT 41.210 25.670 41.440 26.250 ;
        RECT 41.210 24.900 41.440 25.340 ;
        RECT 39.550 23.950 41.440 24.900 ;
        RECT 39.550 22.650 39.900 23.950 ;
        RECT 40.050 23.050 41.050 23.400 ;
        RECT 41.210 23.380 41.440 23.950 ;
        RECT 41.210 22.650 41.440 23.050 ;
        RECT 24.860 21.950 25.090 22.000 ;
        RECT 27.910 21.950 28.140 22.000 ;
        RECT 29.460 21.950 29.690 22.000 ;
        RECT 32.510 21.950 32.740 22.000 ;
        RECT 25.250 21.800 27.750 21.900 ;
        RECT 29.850 21.800 32.350 21.900 ;
        RECT 25.250 21.670 32.350 21.800 ;
        RECT 39.550 21.700 41.440 22.650 ;
        RECT 25.450 21.450 32.100 21.670 ;
        RECT 20.110 21.040 20.340 21.450 ;
        RECT 21.650 21.200 22.600 21.450 ;
        RECT 21.650 21.050 22.980 21.200 ;
        RECT 24.300 21.050 25.300 21.350 ;
        RECT 20.500 20.750 22.980 21.050 ;
        RECT 20.110 20.350 20.340 20.710 ;
        RECT 21.650 20.550 22.980 20.750 ;
        RECT 21.650 20.350 22.600 20.550 ;
        RECT 26.300 20.500 31.550 21.450 ;
        RECT 32.450 21.050 33.450 21.350 ;
        RECT 37.405 21.320 38.295 21.350 ;
        RECT 39.550 21.320 39.900 21.700 ;
        RECT 37.405 20.430 39.900 21.320 ;
        RECT 41.210 21.090 41.440 21.700 ;
        RECT 40.150 21.040 41.050 21.050 ;
        RECT 40.050 20.810 41.050 21.040 ;
        RECT 40.150 20.750 41.050 20.810 ;
        RECT 37.405 20.400 38.295 20.430 ;
        RECT 20.100 19.200 22.600 20.350 ;
        RECT 39.550 20.300 39.900 20.430 ;
        RECT 41.210 20.300 41.440 20.760 ;
        RECT 24.500 20.010 26.460 20.240 ;
        RECT 26.790 20.010 28.750 20.240 ;
        RECT 29.080 20.010 31.040 20.240 ;
        RECT 31.370 20.010 33.330 20.240 ;
        RECT 24.220 19.800 24.450 19.850 ;
        RECT 20.110 18.750 20.340 19.200 ;
        RECT 21.650 18.750 22.600 19.200 ;
        RECT 24.100 18.900 24.500 19.800 ;
        RECT 24.220 18.850 24.450 18.900 ;
        RECT 21.700 18.700 22.600 18.750 ;
        RECT 24.950 18.700 25.850 20.010 ;
        RECT 26.510 19.700 26.740 19.850 ;
        RECT 26.400 19.000 26.850 19.700 ;
        RECT 26.510 18.850 26.740 19.000 ;
        RECT 27.350 18.700 28.250 20.010 ;
        RECT 28.800 19.700 29.030 19.850 ;
        RECT 28.700 19.000 29.150 19.700 ;
        RECT 28.800 18.850 29.030 19.000 ;
        RECT 29.650 18.700 30.550 20.010 ;
        RECT 31.090 19.700 31.320 19.850 ;
        RECT 31.000 19.000 31.450 19.700 ;
        RECT 31.090 18.850 31.320 19.000 ;
        RECT 31.900 18.700 32.800 20.010 ;
        RECT 33.380 19.800 33.610 19.850 ;
        RECT 33.300 18.900 33.700 19.800 ;
        RECT 33.380 18.850 33.610 18.900 ;
        RECT 20.500 18.350 21.500 18.700 ;
        RECT 21.700 18.690 33.300 18.700 ;
        RECT 21.700 18.460 33.330 18.690 ;
        RECT 21.700 18.400 33.300 18.460 ;
        RECT 33.900 18.200 35.250 20.250 ;
        RECT 37.700 18.200 39.400 19.700 ;
        RECT 39.550 19.350 41.500 20.300 ;
        RECT 41.750 19.700 42.500 32.650 ;
        RECT 39.550 18.850 39.900 19.350 ;
        RECT 39.660 18.800 39.890 18.850 ;
        RECT 41.210 18.800 41.440 19.350 ;
        RECT 40.050 18.450 41.050 18.800 ;
        RECT 41.650 18.200 42.500 19.700 ;
        RECT 18.300 17.550 42.500 18.200 ;
        RECT 18.300 16.550 19.350 17.550 ;
        RECT 20.350 16.550 42.500 17.550 ;
        RECT 18.300 15.850 42.500 16.550 ;
      LAYER via ;
        RECT 31.500 38.250 32.500 38.550 ;
        RECT 23.050 36.250 23.900 36.600 ;
        RECT 22.950 35.950 23.900 36.250 ;
        RECT 18.450 18.300 19.250 28.100 ;
        RECT 20.550 27.600 21.450 27.950 ;
        RECT 23.050 31.650 23.900 35.950 ;
        RECT 22.950 31.350 23.900 31.650 ;
        RECT 23.050 27.100 23.900 31.350 ;
        RECT 22.950 26.800 23.900 27.100 ;
        RECT 23.050 26.650 23.900 26.800 ;
        RECT 25.200 35.950 26.100 36.250 ;
        RECT 25.200 31.350 26.100 31.650 ;
        RECT 25.200 26.800 26.100 27.100 ;
        RECT 31.600 35.950 32.500 36.250 ;
        RECT 31.500 33.650 32.500 33.950 ;
        RECT 31.600 31.350 32.500 31.650 ;
        RECT 31.500 29.050 32.500 29.350 ;
        RECT 31.600 26.800 32.500 27.100 ;
        RECT 33.800 36.300 34.650 39.000 ;
        RECT 36.100 38.500 37.050 38.800 ;
        RECT 33.800 36.000 34.750 36.300 ;
        RECT 33.800 31.750 34.650 36.000 ;
        RECT 33.800 31.450 34.750 31.750 ;
        RECT 33.800 29.350 34.650 31.450 ;
        RECT 33.800 28.950 34.700 29.350 ;
        RECT 33.800 27.800 34.650 28.950 ;
        RECT 33.800 27.400 34.700 27.800 ;
        RECT 33.800 27.150 34.650 27.400 ;
        RECT 33.800 26.850 34.750 27.150 ;
        RECT 33.800 26.650 34.650 26.850 ;
        RECT 20.550 23.000 21.450 23.350 ;
        RECT 31.500 24.450 32.500 24.750 ;
        RECT 31.775 24.200 32.325 24.450 ;
        RECT 31.550 22.850 32.400 23.500 ;
        RECT 33.800 23.200 34.700 26.650 ;
        RECT 33.800 22.850 35.050 23.200 ;
        RECT 33.900 22.800 35.050 22.850 ;
        RECT 36.150 37.700 37.100 38.000 ;
        RECT 36.100 36.900 37.050 37.200 ;
        RECT 36.150 36.100 37.100 36.400 ;
        RECT 36.100 35.350 37.050 35.650 ;
        RECT 36.150 34.550 37.100 34.850 ;
        RECT 36.100 33.750 37.050 34.050 ;
        RECT 36.150 32.950 37.100 33.250 ;
        RECT 36.100 32.150 37.050 32.450 ;
        RECT 36.150 31.350 37.100 31.650 ;
        RECT 36.100 30.600 37.050 30.900 ;
        RECT 36.150 29.800 37.100 30.100 ;
        RECT 36.100 29.000 37.050 29.300 ;
        RECT 36.150 28.250 37.100 28.550 ;
        RECT 36.100 27.450 37.050 27.750 ;
        RECT 36.150 26.650 37.100 26.950 ;
        RECT 36.100 25.850 37.050 26.150 ;
        RECT 35.600 25.000 35.900 25.400 ;
        RECT 36.150 25.050 37.100 25.350 ;
        RECT 36.100 24.250 37.050 24.550 ;
        RECT 36.150 23.500 37.100 23.800 ;
        RECT 36.100 22.700 37.050 23.000 ;
        RECT 24.800 22.000 25.100 22.350 ;
        RECT 27.900 22.000 28.200 22.350 ;
        RECT 29.400 22.000 29.700 22.350 ;
        RECT 32.500 22.000 32.800 22.350 ;
        RECT 38.250 22.000 38.850 37.850 ;
        RECT 41.950 35.150 42.350 37.850 ;
        RECT 40.050 34.650 41.000 34.950 ;
        RECT 40.200 34.550 40.950 34.650 ;
        RECT 40.100 32.250 41.000 32.550 ;
        RECT 40.100 29.950 41.000 30.250 ;
        RECT 40.100 27.650 41.000 27.950 ;
        RECT 40.100 25.350 41.000 25.700 ;
        RECT 40.100 23.050 41.000 23.400 ;
        RECT 22.300 20.550 22.950 21.200 ;
        RECT 24.350 21.050 25.250 21.350 ;
        RECT 26.450 20.800 26.850 21.500 ;
        RECT 31.000 20.800 31.400 21.500 ;
        RECT 32.500 21.050 33.400 21.350 ;
        RECT 40.200 20.750 41.000 21.050 ;
        RECT 24.150 18.900 24.450 19.800 ;
        RECT 26.450 19.000 26.800 19.700 ;
        RECT 28.750 19.000 29.100 19.700 ;
        RECT 31.050 19.000 31.400 19.700 ;
        RECT 33.350 18.900 33.650 19.800 ;
        RECT 20.550 18.350 21.450 18.700 ;
        RECT 41.900 20.000 42.300 32.500 ;
        RECT 40.100 18.450 41.000 18.800 ;
        RECT 24.000 17.650 24.500 17.750 ;
        RECT 28.750 17.650 29.100 17.750 ;
        RECT 33.150 17.650 33.650 17.750 ;
        RECT 24.000 17.300 33.650 17.650 ;
        RECT 24.000 17.000 33.600 17.300 ;
      LAYER met2 ;
        RECT 33.800 38.850 34.650 39.050 ;
        RECT 27.910 38.800 29.690 38.840 ;
        RECT 27.900 38.550 32.550 38.800 ;
        RECT 27.910 38.300 32.550 38.550 ;
        RECT 33.800 38.450 37.100 38.850 ;
        RECT 27.910 38.210 32.500 38.300 ;
        RECT 23.050 36.300 23.900 36.650 ;
        RECT 22.950 36.250 23.900 36.300 ;
        RECT 25.200 36.250 26.100 36.300 ;
        RECT 22.900 35.950 26.350 36.250 ;
        RECT 22.950 35.900 23.900 35.950 ;
        RECT 25.200 35.900 26.100 35.950 ;
        RECT 23.050 31.700 23.900 35.900 ;
        RECT 27.910 33.990 29.690 38.210 ;
        RECT 31.500 38.200 32.500 38.210 ;
        RECT 33.800 37.250 34.650 38.450 ;
        RECT 36.100 37.650 42.500 38.050 ;
        RECT 33.800 36.850 37.100 37.250 ;
        RECT 33.800 36.350 34.650 36.850 ;
        RECT 37.900 36.500 42.500 37.650 ;
        RECT 33.800 36.300 34.750 36.350 ;
        RECT 31.600 35.950 34.750 36.300 ;
        RECT 36.100 36.100 42.500 36.500 ;
        RECT 36.150 36.050 37.100 36.100 ;
        RECT 31.600 35.900 32.500 35.950 ;
        RECT 33.800 35.700 34.650 35.950 ;
        RECT 33.800 35.300 37.100 35.700 ;
        RECT 33.800 34.100 34.650 35.300 ;
        RECT 37.900 34.900 42.500 36.100 ;
        RECT 36.100 34.850 42.500 34.900 ;
        RECT 36.100 34.500 41.200 34.850 ;
        RECT 37.900 34.400 41.200 34.500 ;
        RECT 31.500 33.990 32.500 34.000 ;
        RECT 27.910 33.610 32.690 33.990 ;
        RECT 33.800 33.700 37.100 34.100 ;
        RECT 22.950 31.650 23.900 31.700 ;
        RECT 25.200 31.650 26.100 31.700 ;
        RECT 22.900 31.350 26.350 31.650 ;
        RECT 22.950 31.300 23.900 31.350 ;
        RECT 25.200 31.300 26.100 31.350 ;
        RECT 18.450 28.100 19.250 28.150 ;
        RECT 18.450 27.450 21.600 28.100 ;
        RECT 18.450 23.550 19.250 27.450 ;
        RECT 23.050 27.150 23.900 31.300 ;
        RECT 27.910 29.390 29.690 33.610 ;
        RECT 31.500 33.600 32.500 33.610 ;
        RECT 33.800 32.500 34.650 33.700 ;
        RECT 37.900 33.300 39.200 34.400 ;
        RECT 36.100 32.900 39.200 33.300 ;
        RECT 33.800 32.100 37.050 32.500 ;
        RECT 33.800 31.800 34.650 32.100 ;
        RECT 33.800 31.750 34.750 31.800 ;
        RECT 37.900 31.750 39.200 32.900 ;
        RECT 40.050 32.100 42.500 32.650 ;
        RECT 31.600 31.400 34.750 31.750 ;
        RECT 31.600 31.350 34.650 31.400 ;
        RECT 36.100 31.350 39.200 31.750 ;
        RECT 31.600 31.300 32.500 31.350 ;
        RECT 33.800 30.950 34.650 31.350 ;
        RECT 36.150 31.300 37.100 31.350 ;
        RECT 33.800 30.550 37.050 30.950 ;
        RECT 31.500 29.390 32.500 29.400 ;
        RECT 27.910 29.010 32.500 29.390 ;
        RECT 22.950 27.100 23.900 27.150 ;
        RECT 25.200 27.100 26.100 27.150 ;
        RECT 22.900 26.800 26.350 27.100 ;
        RECT 22.950 26.750 23.900 26.800 ;
        RECT 25.200 26.750 26.100 26.800 ;
        RECT 23.050 26.600 23.900 26.750 ;
        RECT 27.910 25.510 29.690 29.010 ;
        RECT 31.500 29.000 32.500 29.010 ;
        RECT 33.800 29.350 34.650 30.550 ;
        RECT 37.900 30.350 39.200 31.350 ;
        RECT 37.900 30.150 41.200 30.350 ;
        RECT 36.100 29.800 41.200 30.150 ;
        RECT 36.100 29.750 39.200 29.800 ;
        RECT 33.800 28.950 37.100 29.350 ;
        RECT 33.800 27.800 34.650 28.950 ;
        RECT 37.900 28.600 39.200 29.750 ;
        RECT 36.100 28.200 39.200 28.600 ;
        RECT 33.800 27.400 37.100 27.800 ;
        RECT 33.800 27.200 34.650 27.400 ;
        RECT 33.800 27.150 34.750 27.200 ;
        RECT 31.600 26.800 34.750 27.150 ;
        RECT 37.900 27.000 39.200 28.200 ;
        RECT 41.750 28.100 42.500 32.100 ;
        RECT 40.050 27.550 42.500 28.100 ;
        RECT 31.600 26.750 32.500 26.800 ;
        RECT 33.800 26.200 34.700 26.800 ;
        RECT 36.100 26.600 39.200 27.000 ;
        RECT 33.800 25.800 37.100 26.200 ;
        RECT 27.920 24.270 29.680 25.510 ;
        RECT 31.775 24.800 32.325 25.370 ;
        RECT 18.450 22.900 21.600 23.550 ;
        RECT 31.500 23.250 32.500 24.800 ;
        RECT 33.800 24.600 34.700 25.800 ;
        RECT 37.900 25.750 39.200 26.600 ;
        RECT 34.900 24.950 35.900 25.450 ;
        RECT 37.900 25.400 41.200 25.750 ;
        RECT 36.100 25.200 41.200 25.400 ;
        RECT 36.100 25.000 39.200 25.200 ;
        RECT 34.900 24.900 35.600 24.950 ;
        RECT 33.800 24.200 37.050 24.600 ;
        RECT 33.800 23.250 34.700 24.200 ;
        RECT 37.900 23.850 39.200 25.000 ;
        RECT 36.100 23.450 39.200 23.850 ;
        RECT 41.750 23.500 42.500 27.550 ;
        RECT 18.450 18.950 19.250 22.900 ;
        RECT 31.550 22.800 32.400 23.250 ;
        RECT 33.800 23.100 35.050 23.250 ;
        RECT 33.800 22.800 37.050 23.100 ;
        RECT 35.150 22.700 37.050 22.800 ;
        RECT 36.100 22.650 37.050 22.700 ;
        RECT 37.900 22.600 39.200 23.450 ;
        RECT 40.050 22.950 42.500 23.500 ;
        RECT 23.500 22.460 24.200 22.500 ;
        RECT 23.475 22.430 24.200 22.460 ;
        RECT 33.525 22.430 34.075 22.460 ;
        RECT 23.475 22.400 28.175 22.430 ;
        RECT 29.425 22.400 34.075 22.430 ;
        RECT 23.475 21.950 28.200 22.400 ;
        RECT 29.400 21.950 34.075 22.400 ;
        RECT 37.900 22.000 41.000 22.600 ;
        RECT 23.475 21.875 28.175 21.950 ;
        RECT 29.425 21.880 34.075 21.950 ;
        RECT 23.475 21.845 24.200 21.875 ;
        RECT 33.525 21.850 34.075 21.880 ;
        RECT 23.500 21.800 24.200 21.845 ;
        RECT 22.300 21.200 22.950 21.230 ;
        RECT 22.300 20.550 23.670 21.200 ;
        RECT 23.950 20.950 25.300 21.400 ;
        RECT 22.300 20.520 22.950 20.550 ;
        RECT 18.450 18.300 21.600 18.950 ;
        RECT 18.450 18.250 19.250 18.300 ;
        RECT 23.950 17.750 24.600 20.950 ;
        RECT 26.350 18.850 26.950 21.600 ;
        RECT 28.650 17.750 29.200 19.850 ;
        RECT 30.900 18.850 31.500 21.600 ;
        RECT 32.400 20.950 33.750 21.400 ;
        RECT 36.385 21.320 37.225 21.495 ;
        RECT 33.100 17.750 33.750 20.950 ;
        RECT 36.360 20.430 38.325 21.320 ;
        RECT 40.200 20.700 41.000 22.000 ;
        RECT 36.385 20.255 37.225 20.430 ;
        RECT 41.750 18.950 42.500 22.950 ;
        RECT 40.050 18.400 42.500 18.950 ;
        RECT 23.950 16.850 33.750 17.750 ;
      LAYER via2 ;
        RECT 28.150 24.750 29.600 25.550 ;
        RECT 31.775 24.775 32.325 25.325 ;
        RECT 22.975 20.550 23.625 21.200 ;
        RECT 36.385 20.300 37.225 21.450 ;
      LAYER met3 ;
        RECT 28.050 25.565 35.000 25.600 ;
        RECT 28.050 25.375 35.565 25.565 ;
        RECT 28.050 24.925 35.600 25.375 ;
        RECT 28.050 24.740 35.565 24.925 ;
        RECT 28.050 24.650 35.000 24.740 ;
        RECT 30.350 24.150 33.200 24.650 ;
        RECT 22.700 20.275 37.250 21.475 ;
  END
END p3_opamp
END LIBRARY

